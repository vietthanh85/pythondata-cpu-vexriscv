// Generator : SpinalHDL v1.7.1    git head : 0444bb76ab1d6e19f0ec46bc03c4769776deb7d5
// Component : VexRiscv
// Git hash  : 11ac8e1c0c66fa0537053980b47757d97dbddf84

`timescale 1ns/1ps

module VexRiscv (
  input      [31:0]   externalResetVector,
  input               timerInterrupt,
  input               softwareInterrupt,
  input      [31:0]   externalInterruptArray,
  output reg          iBusWishbone_CYC,
  output reg          iBusWishbone_STB,
  input               iBusWishbone_ACK,
  output              iBusWishbone_WE,
  output     [29:0]   iBusWishbone_ADR,
  input      [31:0]   iBusWishbone_DAT_MISO,
  output     [31:0]   iBusWishbone_DAT_MOSI,
  output     [3:0]    iBusWishbone_SEL,
  input               iBusWishbone_ERR,
  output     [2:0]    iBusWishbone_CTI,
  output     [1:0]    iBusWishbone_BTE,
  output              dBusWishbone_CYC,
  output              dBusWishbone_STB,
  input               dBusWishbone_ACK,
  output              dBusWishbone_WE,
  output     [29:0]   dBusWishbone_ADR,
  input      [31:0]   dBusWishbone_DAT_MISO,
  output     [31:0]   dBusWishbone_DAT_MOSI,
  output     [3:0]    dBusWishbone_SEL,
  input               dBusWishbone_ERR,
  output     [2:0]    dBusWishbone_CTI,
  output     [1:0]    dBusWishbone_BTE,
  input               clk,
  input               reset
);
  localparam ShiftCtrlEnum_DISABLE_1 = 2'd0;
  localparam ShiftCtrlEnum_SLL_1 = 2'd1;
  localparam ShiftCtrlEnum_SRL_1 = 2'd2;
  localparam ShiftCtrlEnum_SRA_1 = 2'd3;
  localparam EnvCtrlEnum_NONE = 2'd0;
  localparam EnvCtrlEnum_XRET = 2'd1;
  localparam EnvCtrlEnum_WFI = 2'd2;
  localparam EnvCtrlEnum_ECALL = 2'd3;
  localparam BranchCtrlEnum_INC = 2'd0;
  localparam BranchCtrlEnum_B = 2'd1;
  localparam BranchCtrlEnum_JAL = 2'd2;
  localparam BranchCtrlEnum_JALR = 2'd3;
  localparam AluBitwiseCtrlEnum_XOR_1 = 2'd0;
  localparam AluBitwiseCtrlEnum_OR_1 = 2'd1;
  localparam AluBitwiseCtrlEnum_AND_1 = 2'd2;
  localparam Src2CtrlEnum_RS = 2'd0;
  localparam Src2CtrlEnum_IMI = 2'd1;
  localparam Src2CtrlEnum_IMS = 2'd2;
  localparam Src2CtrlEnum_PC = 2'd3;
  localparam AluCtrlEnum_ADD_SUB = 2'd0;
  localparam AluCtrlEnum_SLT_SLTU = 2'd1;
  localparam AluCtrlEnum_BITWISE = 2'd2;
  localparam Src1CtrlEnum_RS = 2'd0;
  localparam Src1CtrlEnum_IMU = 2'd1;
  localparam Src1CtrlEnum_PC_INCREMENT = 2'd2;
  localparam Src1CtrlEnum_URS1 = 2'd3;
  localparam execute_PmpPlugin_fsm_enumDef_BOOT = 3'd0;
  localparam execute_PmpPlugin_fsm_enumDef_stateIdle = 3'd1;
  localparam execute_PmpPlugin_fsm_enumDef_stateWrite = 3'd2;
  localparam execute_PmpPlugin_fsm_enumDef_stateCfg = 3'd3;
  localparam execute_PmpPlugin_fsm_enumDef_stateAddr = 3'd4;

  reg        [31:0]   PmpPlugin_setter_io_addr;
  wire                IBusCachedPlugin_cache_io_flush;
  wire                IBusCachedPlugin_cache_io_cpu_prefetch_isValid;
  wire                IBusCachedPlugin_cache_io_cpu_fetch_isValid;
  wire                IBusCachedPlugin_cache_io_cpu_fetch_isStuck;
  wire                IBusCachedPlugin_cache_io_cpu_fetch_isRemoved;
  wire                IBusCachedPlugin_cache_io_cpu_decode_isValid;
  wire                IBusCachedPlugin_cache_io_cpu_decode_isStuck;
  wire                IBusCachedPlugin_cache_io_cpu_decode_isUser;
  reg                 IBusCachedPlugin_cache_io_cpu_fill_valid;
  wire                dataCache_1_io_cpu_execute_isValid;
  wire       [31:0]   dataCache_1_io_cpu_execute_address;
  wire                dataCache_1_io_cpu_memory_isValid;
  wire       [31:0]   dataCache_1_io_cpu_memory_address;
  reg                 dataCache_1_io_cpu_memory_mmuRsp_isIoAccess;
  reg                 dataCache_1_io_cpu_writeBack_isValid;
  wire                dataCache_1_io_cpu_writeBack_isUser;
  wire       [31:0]   dataCache_1_io_cpu_writeBack_storeData;
  wire       [31:0]   dataCache_1_io_cpu_writeBack_address;
  wire                dataCache_1_io_cpu_writeBack_fence_SW;
  wire                dataCache_1_io_cpu_writeBack_fence_SR;
  wire                dataCache_1_io_cpu_writeBack_fence_SO;
  wire                dataCache_1_io_cpu_writeBack_fence_SI;
  wire                dataCache_1_io_cpu_writeBack_fence_PW;
  wire                dataCache_1_io_cpu_writeBack_fence_PR;
  wire                dataCache_1_io_cpu_writeBack_fence_PO;
  wire                dataCache_1_io_cpu_writeBack_fence_PI;
  wire       [3:0]    dataCache_1_io_cpu_writeBack_fence_FM;
  wire                dataCache_1_io_cpu_flush_valid;
  wire                dataCache_1_io_cpu_flush_payload_singleLine;
  wire       [6:0]    dataCache_1_io_cpu_flush_payload_lineId;
  wire                dataCache_1_io_mem_cmd_ready;
  wire       [31:0]   _zz_PmpPlugin_pmpaddr_port0;
  wire       [31:0]   _zz_PmpPlugin_pmpaddr_port2;
  reg        [31:0]   _zz_RegFilePlugin_regFile_port0;
  reg        [31:0]   _zz_RegFilePlugin_regFile_port1;
  wire       [24:0]   PmpPlugin_setter_io_base;
  wire       [24:0]   PmpPlugin_setter_io_mask;
  wire                IBusCachedPlugin_cache_io_cpu_prefetch_haltIt;
  wire       [31:0]   IBusCachedPlugin_cache_io_cpu_fetch_data;
  wire       [31:0]   IBusCachedPlugin_cache_io_cpu_fetch_physicalAddress;
  wire                IBusCachedPlugin_cache_io_cpu_decode_error;
  wire                IBusCachedPlugin_cache_io_cpu_decode_mmuRefilling;
  wire                IBusCachedPlugin_cache_io_cpu_decode_mmuException;
  wire       [31:0]   IBusCachedPlugin_cache_io_cpu_decode_data;
  wire                IBusCachedPlugin_cache_io_cpu_decode_cacheMiss;
  wire       [31:0]   IBusCachedPlugin_cache_io_cpu_decode_physicalAddress;
  wire                IBusCachedPlugin_cache_io_mem_cmd_valid;
  wire       [31:0]   IBusCachedPlugin_cache_io_mem_cmd_payload_address;
  wire       [2:0]    IBusCachedPlugin_cache_io_mem_cmd_payload_size;
  wire                dataCache_1_io_cpu_execute_haltIt;
  wire                dataCache_1_io_cpu_execute_refilling;
  wire                dataCache_1_io_cpu_memory_isWrite;
  wire                dataCache_1_io_cpu_writeBack_haltIt;
  wire       [31:0]   dataCache_1_io_cpu_writeBack_data;
  wire                dataCache_1_io_cpu_writeBack_mmuException;
  wire                dataCache_1_io_cpu_writeBack_unalignedAccess;
  wire                dataCache_1_io_cpu_writeBack_accessError;
  wire                dataCache_1_io_cpu_writeBack_isWrite;
  wire                dataCache_1_io_cpu_writeBack_keepMemRspData;
  wire                dataCache_1_io_cpu_writeBack_exclusiveOk;
  wire                dataCache_1_io_cpu_flush_ready;
  wire                dataCache_1_io_cpu_redo;
  wire                dataCache_1_io_mem_cmd_valid;
  wire                dataCache_1_io_mem_cmd_payload_wr;
  wire                dataCache_1_io_mem_cmd_payload_uncached;
  wire       [31:0]   dataCache_1_io_mem_cmd_payload_address;
  wire       [31:0]   dataCache_1_io_mem_cmd_payload_data;
  wire       [3:0]    dataCache_1_io_mem_cmd_payload_mask;
  wire       [2:0]    dataCache_1_io_mem_cmd_payload_size;
  wire                dataCache_1_io_mem_cmd_payload_last;
  wire       [51:0]   _zz_memory_MUL_LOW;
  wire       [51:0]   _zz_memory_MUL_LOW_1;
  wire       [51:0]   _zz_memory_MUL_LOW_2;
  wire       [51:0]   _zz_memory_MUL_LOW_3;
  wire       [32:0]   _zz_memory_MUL_LOW_4;
  wire       [51:0]   _zz_memory_MUL_LOW_5;
  wire       [49:0]   _zz_memory_MUL_LOW_6;
  wire       [51:0]   _zz_memory_MUL_LOW_7;
  wire       [49:0]   _zz_memory_MUL_LOW_8;
  wire       [31:0]   _zz_execute_SHIFT_RIGHT;
  wire       [32:0]   _zz_execute_SHIFT_RIGHT_1;
  wire       [32:0]   _zz_execute_SHIFT_RIGHT_2;
  wire       [31:0]   _zz_decode_LEGAL_INSTRUCTION;
  wire       [31:0]   _zz_decode_LEGAL_INSTRUCTION_1;
  wire       [31:0]   _zz_decode_LEGAL_INSTRUCTION_2;
  wire                _zz_decode_LEGAL_INSTRUCTION_3;
  wire       [0:0]    _zz_decode_LEGAL_INSTRUCTION_4;
  wire       [13:0]   _zz_decode_LEGAL_INSTRUCTION_5;
  wire       [31:0]   _zz_decode_LEGAL_INSTRUCTION_6;
  wire       [31:0]   _zz_decode_LEGAL_INSTRUCTION_7;
  wire       [31:0]   _zz_decode_LEGAL_INSTRUCTION_8;
  wire                _zz_decode_LEGAL_INSTRUCTION_9;
  wire       [0:0]    _zz_decode_LEGAL_INSTRUCTION_10;
  wire       [7:0]    _zz_decode_LEGAL_INSTRUCTION_11;
  wire       [31:0]   _zz_decode_LEGAL_INSTRUCTION_12;
  wire       [31:0]   _zz_decode_LEGAL_INSTRUCTION_13;
  wire       [31:0]   _zz_decode_LEGAL_INSTRUCTION_14;
  wire                _zz_decode_LEGAL_INSTRUCTION_15;
  wire       [0:0]    _zz_decode_LEGAL_INSTRUCTION_16;
  wire       [1:0]    _zz_decode_LEGAL_INSTRUCTION_17;
  wire       [3:0]    _zz__zz_IBusCachedPlugin_jump_pcLoad_payload_1;
  reg        [31:0]   _zz_IBusCachedPlugin_jump_pcLoad_payload_5;
  wire       [1:0]    _zz_IBusCachedPlugin_jump_pcLoad_payload_6;
  wire       [31:0]   _zz_IBusCachedPlugin_fetchPc_pc;
  wire       [2:0]    _zz_IBusCachedPlugin_fetchPc_pc_1;
  wire       [11:0]   _zz__zz_IBusCachedPlugin_decodePrediction_cmd_hadBranch;
  wire       [31:0]   _zz_IBusCachedPlugin_decodePrediction_cmd_hadBranch_2;
  wire       [19:0]   _zz__zz_3;
  wire       [11:0]   _zz__zz_5;
  wire       [31:0]   _zz__zz_7;
  wire       [31:0]   _zz__zz_7_1;
  wire       [19:0]   _zz__zz_IBusCachedPlugin_predictionJumpInterface_payload;
  wire       [11:0]   _zz__zz_IBusCachedPlugin_predictionJumpInterface_payload_2;
  wire                _zz_IBusCachedPlugin_predictionJumpInterface_payload_4;
  wire                _zz_IBusCachedPlugin_predictionJumpInterface_payload_5;
  wire                _zz_IBusCachedPlugin_predictionJumpInterface_payload_6;
  wire       [26:0]   _zz_io_cpu_flush_payload_lineId;
  wire       [26:0]   _zz_io_cpu_flush_payload_lineId_1;
  wire       [2:0]    _zz_DBusCachedPlugin_exceptionBus_payload_code;
  wire       [2:0]    _zz_DBusCachedPlugin_exceptionBus_payload_code_1;
  reg        [7:0]    _zz_writeBack_DBusCachedPlugin_rspShifted;
  wire       [1:0]    _zz_writeBack_DBusCachedPlugin_rspShifted_1;
  reg        [7:0]    _zz_writeBack_DBusCachedPlugin_rspShifted_2;
  wire       [0:0]    _zz_writeBack_DBusCachedPlugin_rspShifted_3;
  reg        [7:0]    _zz_when_PmpPlugin_l246;
  reg        [24:0]   _zz_PmpPlugin_dGuard_hits_0_1;
  wire       [3:0]    _zz_PmpPlugin_dGuard_hits_0_2;
  reg        [24:0]   _zz_PmpPlugin_dGuard_hits_0_3;
  wire       [3:0]    _zz_PmpPlugin_dGuard_hits_0_4;
  reg        [24:0]   _zz_PmpPlugin_dGuard_hits_1;
  wire       [3:0]    _zz_PmpPlugin_dGuard_hits_1_1;
  reg        [24:0]   _zz_PmpPlugin_dGuard_hits_1_2;
  wire       [3:0]    _zz_PmpPlugin_dGuard_hits_1_3;
  reg        [24:0]   _zz_PmpPlugin_dGuard_hits_2;
  wire       [3:0]    _zz_PmpPlugin_dGuard_hits_2_1;
  reg        [24:0]   _zz_PmpPlugin_dGuard_hits_2_2;
  wire       [3:0]    _zz_PmpPlugin_dGuard_hits_2_3;
  reg        [24:0]   _zz_PmpPlugin_dGuard_hits_3;
  wire       [3:0]    _zz_PmpPlugin_dGuard_hits_3_1;
  reg        [24:0]   _zz_PmpPlugin_dGuard_hits_3_2;
  wire       [3:0]    _zz_PmpPlugin_dGuard_hits_3_3;
  reg        [24:0]   _zz_PmpPlugin_dGuard_hits_4;
  wire       [3:0]    _zz_PmpPlugin_dGuard_hits_4_1;
  reg        [24:0]   _zz_PmpPlugin_dGuard_hits_4_2;
  wire       [3:0]    _zz_PmpPlugin_dGuard_hits_4_3;
  reg        [24:0]   _zz_PmpPlugin_dGuard_hits_5;
  wire       [3:0]    _zz_PmpPlugin_dGuard_hits_5_1;
  reg        [24:0]   _zz_PmpPlugin_dGuard_hits_5_2;
  wire       [3:0]    _zz_PmpPlugin_dGuard_hits_5_3;
  reg        [24:0]   _zz_PmpPlugin_dGuard_hits_6;
  wire       [3:0]    _zz_PmpPlugin_dGuard_hits_6_1;
  reg        [24:0]   _zz_PmpPlugin_dGuard_hits_6_2;
  wire       [3:0]    _zz_PmpPlugin_dGuard_hits_6_3;
  reg        [24:0]   _zz_PmpPlugin_dGuard_hits_7;
  wire       [3:0]    _zz_PmpPlugin_dGuard_hits_7_1;
  reg        [24:0]   _zz_PmpPlugin_dGuard_hits_7_2;
  wire       [3:0]    _zz_PmpPlugin_dGuard_hits_7_3;
  reg        [24:0]   _zz_PmpPlugin_dGuard_hits_8;
  wire       [3:0]    _zz_PmpPlugin_dGuard_hits_8_1;
  reg        [24:0]   _zz_PmpPlugin_dGuard_hits_8_2;
  wire       [3:0]    _zz_PmpPlugin_dGuard_hits_8_3;
  reg        [24:0]   _zz_PmpPlugin_dGuard_hits_9;
  wire       [3:0]    _zz_PmpPlugin_dGuard_hits_9_1;
  reg        [24:0]   _zz_PmpPlugin_dGuard_hits_9_2;
  wire       [3:0]    _zz_PmpPlugin_dGuard_hits_9_3;
  reg        [24:0]   _zz_PmpPlugin_dGuard_hits_10;
  wire       [3:0]    _zz_PmpPlugin_dGuard_hits_10_1;
  reg        [24:0]   _zz_PmpPlugin_dGuard_hits_10_2;
  wire       [3:0]    _zz_PmpPlugin_dGuard_hits_10_3;
  reg        [24:0]   _zz_PmpPlugin_dGuard_hits_11;
  wire       [3:0]    _zz_PmpPlugin_dGuard_hits_11_1;
  reg        [24:0]   _zz_PmpPlugin_dGuard_hits_11_2;
  wire       [3:0]    _zz_PmpPlugin_dGuard_hits_11_3;
  reg        [24:0]   _zz_PmpPlugin_dGuard_hits_12;
  wire       [3:0]    _zz_PmpPlugin_dGuard_hits_12_1;
  reg        [24:0]   _zz_PmpPlugin_dGuard_hits_12_2;
  wire       [3:0]    _zz_PmpPlugin_dGuard_hits_12_3;
  reg        [24:0]   _zz_PmpPlugin_dGuard_hits_13;
  wire       [3:0]    _zz_PmpPlugin_dGuard_hits_13_1;
  reg        [24:0]   _zz_PmpPlugin_dGuard_hits_13_2;
  wire       [3:0]    _zz_PmpPlugin_dGuard_hits_13_3;
  reg        [24:0]   _zz_PmpPlugin_dGuard_hits_14;
  wire       [3:0]    _zz_PmpPlugin_dGuard_hits_14_1;
  reg        [24:0]   _zz_PmpPlugin_dGuard_hits_14_2;
  wire       [3:0]    _zz_PmpPlugin_dGuard_hits_14_3;
  reg        [24:0]   _zz_PmpPlugin_dGuard_hits_15;
  wire       [3:0]    _zz_PmpPlugin_dGuard_hits_15_1;
  reg        [24:0]   _zz_PmpPlugin_dGuard_hits_15_2;
  wire       [3:0]    _zz_PmpPlugin_dGuard_hits_15_3;
  wire       [0:0]    _zz_when_PmpPlugin_l277;
  wire       [5:0]    _zz_when_PmpPlugin_l277_1;
  wire       [0:0]    _zz__zz_DBusCachedPlugin_mmuBus_rsp_allowRead;
  wire       [4:0]    _zz__zz_DBusCachedPlugin_mmuBus_rsp_allowRead_1;
  wire       [15:0]   _zz__zz_DBusCachedPlugin_mmuBus_rsp_allowRead_1_1;
  reg                 _zz_DBusCachedPlugin_mmuBus_rsp_allowRead_17;
  wire       [3:0]    _zz_DBusCachedPlugin_mmuBus_rsp_allowRead_18;
  wire       [0:0]    _zz__zz_DBusCachedPlugin_mmuBus_rsp_allowWrite;
  wire       [4:0]    _zz__zz_DBusCachedPlugin_mmuBus_rsp_allowWrite_1;
  wire       [15:0]   _zz__zz_DBusCachedPlugin_mmuBus_rsp_allowWrite_1_1;
  reg                 _zz_DBusCachedPlugin_mmuBus_rsp_allowWrite_17;
  wire       [3:0]    _zz_DBusCachedPlugin_mmuBus_rsp_allowWrite_18;
  reg        [24:0]   _zz_PmpPlugin_iGuard_hits_0_1;
  wire       [3:0]    _zz_PmpPlugin_iGuard_hits_0_2;
  reg        [24:0]   _zz_PmpPlugin_iGuard_hits_0_3;
  wire       [3:0]    _zz_PmpPlugin_iGuard_hits_0_4;
  reg        [24:0]   _zz_PmpPlugin_iGuard_hits_1;
  wire       [3:0]    _zz_PmpPlugin_iGuard_hits_1_1;
  reg        [24:0]   _zz_PmpPlugin_iGuard_hits_1_2;
  wire       [3:0]    _zz_PmpPlugin_iGuard_hits_1_3;
  reg        [24:0]   _zz_PmpPlugin_iGuard_hits_2;
  wire       [3:0]    _zz_PmpPlugin_iGuard_hits_2_1;
  reg        [24:0]   _zz_PmpPlugin_iGuard_hits_2_2;
  wire       [3:0]    _zz_PmpPlugin_iGuard_hits_2_3;
  reg        [24:0]   _zz_PmpPlugin_iGuard_hits_3;
  wire       [3:0]    _zz_PmpPlugin_iGuard_hits_3_1;
  reg        [24:0]   _zz_PmpPlugin_iGuard_hits_3_2;
  wire       [3:0]    _zz_PmpPlugin_iGuard_hits_3_3;
  reg        [24:0]   _zz_PmpPlugin_iGuard_hits_4;
  wire       [3:0]    _zz_PmpPlugin_iGuard_hits_4_1;
  reg        [24:0]   _zz_PmpPlugin_iGuard_hits_4_2;
  wire       [3:0]    _zz_PmpPlugin_iGuard_hits_4_3;
  reg        [24:0]   _zz_PmpPlugin_iGuard_hits_5;
  wire       [3:0]    _zz_PmpPlugin_iGuard_hits_5_1;
  reg        [24:0]   _zz_PmpPlugin_iGuard_hits_5_2;
  wire       [3:0]    _zz_PmpPlugin_iGuard_hits_5_3;
  reg        [24:0]   _zz_PmpPlugin_iGuard_hits_6;
  wire       [3:0]    _zz_PmpPlugin_iGuard_hits_6_1;
  reg        [24:0]   _zz_PmpPlugin_iGuard_hits_6_2;
  wire       [3:0]    _zz_PmpPlugin_iGuard_hits_6_3;
  reg        [24:0]   _zz_PmpPlugin_iGuard_hits_7;
  wire       [3:0]    _zz_PmpPlugin_iGuard_hits_7_1;
  reg        [24:0]   _zz_PmpPlugin_iGuard_hits_7_2;
  wire       [3:0]    _zz_PmpPlugin_iGuard_hits_7_3;
  reg        [24:0]   _zz_PmpPlugin_iGuard_hits_8;
  wire       [3:0]    _zz_PmpPlugin_iGuard_hits_8_1;
  reg        [24:0]   _zz_PmpPlugin_iGuard_hits_8_2;
  wire       [3:0]    _zz_PmpPlugin_iGuard_hits_8_3;
  reg        [24:0]   _zz_PmpPlugin_iGuard_hits_9;
  wire       [3:0]    _zz_PmpPlugin_iGuard_hits_9_1;
  reg        [24:0]   _zz_PmpPlugin_iGuard_hits_9_2;
  wire       [3:0]    _zz_PmpPlugin_iGuard_hits_9_3;
  reg        [24:0]   _zz_PmpPlugin_iGuard_hits_10;
  wire       [3:0]    _zz_PmpPlugin_iGuard_hits_10_1;
  reg        [24:0]   _zz_PmpPlugin_iGuard_hits_10_2;
  wire       [3:0]    _zz_PmpPlugin_iGuard_hits_10_3;
  reg        [24:0]   _zz_PmpPlugin_iGuard_hits_11;
  wire       [3:0]    _zz_PmpPlugin_iGuard_hits_11_1;
  reg        [24:0]   _zz_PmpPlugin_iGuard_hits_11_2;
  wire       [3:0]    _zz_PmpPlugin_iGuard_hits_11_3;
  reg        [24:0]   _zz_PmpPlugin_iGuard_hits_12;
  wire       [3:0]    _zz_PmpPlugin_iGuard_hits_12_1;
  reg        [24:0]   _zz_PmpPlugin_iGuard_hits_12_2;
  wire       [3:0]    _zz_PmpPlugin_iGuard_hits_12_3;
  reg        [24:0]   _zz_PmpPlugin_iGuard_hits_13;
  wire       [3:0]    _zz_PmpPlugin_iGuard_hits_13_1;
  reg        [24:0]   _zz_PmpPlugin_iGuard_hits_13_2;
  wire       [3:0]    _zz_PmpPlugin_iGuard_hits_13_3;
  reg        [24:0]   _zz_PmpPlugin_iGuard_hits_14;
  wire       [3:0]    _zz_PmpPlugin_iGuard_hits_14_1;
  reg        [24:0]   _zz_PmpPlugin_iGuard_hits_14_2;
  wire       [3:0]    _zz_PmpPlugin_iGuard_hits_14_3;
  reg        [24:0]   _zz_PmpPlugin_iGuard_hits_15;
  wire       [3:0]    _zz_PmpPlugin_iGuard_hits_15_1;
  reg        [24:0]   _zz_PmpPlugin_iGuard_hits_15_2;
  wire       [3:0]    _zz_PmpPlugin_iGuard_hits_15_3;
  wire       [0:0]    _zz_when_PmpPlugin_l299;
  wire       [5:0]    _zz_when_PmpPlugin_l299_1;
  wire       [0:0]    _zz__zz_IBusCachedPlugin_mmuBus_rsp_allowExecute;
  wire       [4:0]    _zz__zz_IBusCachedPlugin_mmuBus_rsp_allowExecute_1;
  wire       [15:0]   _zz__zz_IBusCachedPlugin_mmuBus_rsp_allowExecute_1_1;
  reg                 _zz_IBusCachedPlugin_mmuBus_rsp_allowExecute_17;
  wire       [3:0]    _zz_IBusCachedPlugin_mmuBus_rsp_allowExecute_18;
  wire       [31:0]   _zz__zz_decode_IS_RS2_SIGNED;
  wire       [31:0]   _zz__zz_decode_IS_RS2_SIGNED_1;
  wire                _zz__zz_decode_IS_RS2_SIGNED_2;
  wire       [0:0]    _zz__zz_decode_IS_RS2_SIGNED_3;
  wire                _zz__zz_decode_IS_RS2_SIGNED_4;
  wire       [31:0]   _zz__zz_decode_IS_RS2_SIGNED_5;
  wire       [0:0]    _zz__zz_decode_IS_RS2_SIGNED_6;
  wire                _zz__zz_decode_IS_RS2_SIGNED_7;
  wire                _zz__zz_decode_IS_RS2_SIGNED_8;
  wire       [24:0]   _zz__zz_decode_IS_RS2_SIGNED_9;
  wire       [0:0]    _zz__zz_decode_IS_RS2_SIGNED_10;
  wire       [0:0]    _zz__zz_decode_IS_RS2_SIGNED_11;
  wire       [31:0]   _zz__zz_decode_IS_RS2_SIGNED_12;
  wire       [0:0]    _zz__zz_decode_IS_RS2_SIGNED_13;
  wire       [31:0]   _zz__zz_decode_IS_RS2_SIGNED_14;
  wire                _zz__zz_decode_IS_RS2_SIGNED_15;
  wire                _zz__zz_decode_IS_RS2_SIGNED_16;
  wire                _zz__zz_decode_IS_RS2_SIGNED_17;
  wire       [0:0]    _zz__zz_decode_IS_RS2_SIGNED_18;
  wire       [0:0]    _zz__zz_decode_IS_RS2_SIGNED_19;
  wire       [31:0]   _zz__zz_decode_IS_RS2_SIGNED_20;
  wire       [1:0]    _zz__zz_decode_IS_RS2_SIGNED_21;
  wire       [31:0]   _zz__zz_decode_IS_RS2_SIGNED_22;
  wire       [31:0]   _zz__zz_decode_IS_RS2_SIGNED_23;
  wire       [31:0]   _zz__zz_decode_IS_RS2_SIGNED_24;
  wire       [31:0]   _zz__zz_decode_IS_RS2_SIGNED_25;
  wire       [20:0]   _zz__zz_decode_IS_RS2_SIGNED_26;
  wire       [0:0]    _zz__zz_decode_IS_RS2_SIGNED_27;
  wire       [31:0]   _zz__zz_decode_IS_RS2_SIGNED_28;
  wire                _zz__zz_decode_IS_RS2_SIGNED_29;
  wire       [31:0]   _zz__zz_decode_IS_RS2_SIGNED_30;
  wire       [31:0]   _zz__zz_decode_IS_RS2_SIGNED_31;
  wire       [0:0]    _zz__zz_decode_IS_RS2_SIGNED_32;
  wire                _zz__zz_decode_IS_RS2_SIGNED_33;
  wire       [17:0]   _zz__zz_decode_IS_RS2_SIGNED_34;
  wire       [1:0]    _zz__zz_decode_IS_RS2_SIGNED_35;
  wire       [31:0]   _zz__zz_decode_IS_RS2_SIGNED_36;
  wire       [31:0]   _zz__zz_decode_IS_RS2_SIGNED_37;
  wire                _zz__zz_decode_IS_RS2_SIGNED_38;
  wire       [31:0]   _zz__zz_decode_IS_RS2_SIGNED_39;
  wire       [0:0]    _zz__zz_decode_IS_RS2_SIGNED_40;
  wire                _zz__zz_decode_IS_RS2_SIGNED_41;
  wire                _zz__zz_decode_IS_RS2_SIGNED_42;
  wire       [14:0]   _zz__zz_decode_IS_RS2_SIGNED_43;
  wire       [0:0]    _zz__zz_decode_IS_RS2_SIGNED_44;
  wire       [31:0]   _zz__zz_decode_IS_RS2_SIGNED_45;
  wire       [3:0]    _zz__zz_decode_IS_RS2_SIGNED_46;
  wire       [31:0]   _zz__zz_decode_IS_RS2_SIGNED_47;
  wire       [31:0]   _zz__zz_decode_IS_RS2_SIGNED_48;
  wire                _zz__zz_decode_IS_RS2_SIGNED_49;
  wire       [31:0]   _zz__zz_decode_IS_RS2_SIGNED_50;
  wire       [0:0]    _zz__zz_decode_IS_RS2_SIGNED_51;
  wire       [31:0]   _zz__zz_decode_IS_RS2_SIGNED_52;
  wire       [31:0]   _zz__zz_decode_IS_RS2_SIGNED_53;
  wire       [0:0]    _zz__zz_decode_IS_RS2_SIGNED_54;
  wire       [0:0]    _zz__zz_decode_IS_RS2_SIGNED_55;
  wire       [31:0]   _zz__zz_decode_IS_RS2_SIGNED_56;
  wire                _zz__zz_decode_IS_RS2_SIGNED_57;
  wire                _zz__zz_decode_IS_RS2_SIGNED_58;
  wire       [31:0]   _zz__zz_decode_IS_RS2_SIGNED_59;
  wire       [0:0]    _zz__zz_decode_IS_RS2_SIGNED_60;
  wire       [2:0]    _zz__zz_decode_IS_RS2_SIGNED_61;
  wire                _zz__zz_decode_IS_RS2_SIGNED_62;
  wire       [31:0]   _zz__zz_decode_IS_RS2_SIGNED_63;
  wire       [0:0]    _zz__zz_decode_IS_RS2_SIGNED_64;
  wire       [31:0]   _zz__zz_decode_IS_RS2_SIGNED_65;
  wire       [31:0]   _zz__zz_decode_IS_RS2_SIGNED_66;
  wire       [0:0]    _zz__zz_decode_IS_RS2_SIGNED_67;
  wire       [31:0]   _zz__zz_decode_IS_RS2_SIGNED_68;
  wire       [31:0]   _zz__zz_decode_IS_RS2_SIGNED_69;
  wire       [0:0]    _zz__zz_decode_IS_RS2_SIGNED_70;
  wire       [0:0]    _zz__zz_decode_IS_RS2_SIGNED_71;
  wire       [3:0]    _zz__zz_decode_IS_RS2_SIGNED_72;
  wire                _zz__zz_decode_IS_RS2_SIGNED_73;
  wire       [31:0]   _zz__zz_decode_IS_RS2_SIGNED_74;
  wire       [0:0]    _zz__zz_decode_IS_RS2_SIGNED_75;
  wire       [31:0]   _zz__zz_decode_IS_RS2_SIGNED_76;
  wire       [31:0]   _zz__zz_decode_IS_RS2_SIGNED_77;
  wire       [1:0]    _zz__zz_decode_IS_RS2_SIGNED_78;
  wire                _zz__zz_decode_IS_RS2_SIGNED_79;
  wire       [31:0]   _zz__zz_decode_IS_RS2_SIGNED_80;
  wire                _zz__zz_decode_IS_RS2_SIGNED_81;
  wire       [31:0]   _zz__zz_decode_IS_RS2_SIGNED_82;
  wire       [10:0]   _zz__zz_decode_IS_RS2_SIGNED_83;
  wire       [5:0]    _zz__zz_decode_IS_RS2_SIGNED_84;
  wire       [0:0]    _zz__zz_decode_IS_RS2_SIGNED_85;
  wire       [31:0]   _zz__zz_decode_IS_RS2_SIGNED_86;
  wire       [31:0]   _zz__zz_decode_IS_RS2_SIGNED_87;
  wire       [3:0]    _zz__zz_decode_IS_RS2_SIGNED_88;
  wire                _zz__zz_decode_IS_RS2_SIGNED_89;
  wire       [31:0]   _zz__zz_decode_IS_RS2_SIGNED_90;
  wire       [0:0]    _zz__zz_decode_IS_RS2_SIGNED_91;
  wire       [31:0]   _zz__zz_decode_IS_RS2_SIGNED_92;
  wire       [31:0]   _zz__zz_decode_IS_RS2_SIGNED_93;
  wire       [1:0]    _zz__zz_decode_IS_RS2_SIGNED_94;
  wire                _zz__zz_decode_IS_RS2_SIGNED_95;
  wire                _zz__zz_decode_IS_RS2_SIGNED_96;
  wire                _zz__zz_decode_IS_RS2_SIGNED_97;
  wire       [0:0]    _zz__zz_decode_IS_RS2_SIGNED_98;
  wire       [0:0]    _zz__zz_decode_IS_RS2_SIGNED_99;
  wire       [31:0]   _zz__zz_decode_IS_RS2_SIGNED_100;
  wire       [31:0]   _zz__zz_decode_IS_RS2_SIGNED_101;
  wire       [0:0]    _zz__zz_decode_IS_RS2_SIGNED_102;
  wire       [1:0]    _zz__zz_decode_IS_RS2_SIGNED_103;
  wire                _zz__zz_decode_IS_RS2_SIGNED_104;
  wire       [31:0]   _zz__zz_decode_IS_RS2_SIGNED_105;
  wire       [7:0]    _zz__zz_decode_IS_RS2_SIGNED_106;
  wire                _zz__zz_decode_IS_RS2_SIGNED_107;
  wire                _zz__zz_decode_IS_RS2_SIGNED_108;
  wire       [31:0]   _zz__zz_decode_IS_RS2_SIGNED_109;
  wire       [0:0]    _zz__zz_decode_IS_RS2_SIGNED_110;
  wire       [0:0]    _zz__zz_decode_IS_RS2_SIGNED_111;
  wire       [31:0]   _zz__zz_decode_IS_RS2_SIGNED_112;
  wire       [31:0]   _zz__zz_decode_IS_RS2_SIGNED_113;
  wire       [5:0]    _zz__zz_decode_IS_RS2_SIGNED_114;
  wire                _zz__zz_decode_IS_RS2_SIGNED_115;
  wire       [0:0]    _zz__zz_decode_IS_RS2_SIGNED_116;
  wire       [31:0]   _zz__zz_decode_IS_RS2_SIGNED_117;
  wire       [3:0]    _zz__zz_decode_IS_RS2_SIGNED_118;
  wire                _zz__zz_decode_IS_RS2_SIGNED_119;
  wire       [0:0]    _zz__zz_decode_IS_RS2_SIGNED_120;
  wire       [31:0]   _zz__zz_decode_IS_RS2_SIGNED_121;
  wire       [0:0]    _zz__zz_decode_IS_RS2_SIGNED_122;
  wire       [31:0]   _zz__zz_decode_IS_RS2_SIGNED_123;
  wire       [0:0]    _zz__zz_decode_IS_RS2_SIGNED_124;
  wire       [0:0]    _zz__zz_decode_IS_RS2_SIGNED_125;
  wire       [31:0]   _zz__zz_decode_IS_RS2_SIGNED_126;
  wire       [3:0]    _zz__zz_decode_IS_RS2_SIGNED_127;
  wire                _zz__zz_decode_IS_RS2_SIGNED_128;
  wire                _zz__zz_decode_IS_RS2_SIGNED_129;
  wire       [0:0]    _zz__zz_decode_IS_RS2_SIGNED_130;
  wire       [31:0]   _zz__zz_decode_IS_RS2_SIGNED_131;
  wire       [0:0]    _zz__zz_decode_IS_RS2_SIGNED_132;
  wire       [31:0]   _zz__zz_decode_IS_RS2_SIGNED_133;
  wire       [0:0]    _zz__zz_decode_IS_RS2_SIGNED_134;
  wire       [0:0]    _zz__zz_decode_IS_RS2_SIGNED_135;
  wire       [31:0]   _zz__zz_decode_IS_RS2_SIGNED_136;
  wire       [0:0]    _zz__zz_decode_IS_RS2_SIGNED_137;
  wire       [1:0]    _zz__zz_decode_IS_RS2_SIGNED_138;
  wire       [1:0]    _zz__zz_decode_IS_RS2_SIGNED_139;
  wire       [31:0]   _zz__zz_decode_IS_RS2_SIGNED_140;
  wire       [31:0]   _zz__zz_decode_IS_RS2_SIGNED_141;
  wire       [0:0]    _zz__zz_decode_IS_RS2_SIGNED_142;
  wire       [31:0]   _zz__zz_decode_IS_RS2_SIGNED_143;
  wire                _zz_RegFilePlugin_regFile_port;
  wire                _zz_decode_RegFilePlugin_rs1Data;
  wire                _zz_RegFilePlugin_regFile_port_1;
  wire                _zz_decode_RegFilePlugin_rs2Data;
  wire       [0:0]    _zz__zz_execute_REGFILE_WRITE_DATA;
  wire       [2:0]    _zz__zz_execute_SRC1;
  wire       [4:0]    _zz__zz_execute_SRC1_1;
  wire       [11:0]   _zz__zz_execute_SRC2_3;
  wire       [31:0]   _zz_execute_SrcPlugin_addSub;
  wire       [31:0]   _zz_execute_SrcPlugin_addSub_1;
  wire       [31:0]   _zz_execute_SrcPlugin_addSub_2;
  wire       [31:0]   _zz_execute_SrcPlugin_addSub_3;
  wire       [31:0]   _zz_execute_SrcPlugin_addSub_4;
  wire       [31:0]   _zz_execute_SrcPlugin_addSub_5;
  wire       [31:0]   _zz_execute_SrcPlugin_addSub_6;
  wire       [19:0]   _zz__zz_execute_BranchPlugin_missAlignedTarget_2;
  wire       [11:0]   _zz__zz_execute_BranchPlugin_missAlignedTarget_4;
  wire       [31:0]   _zz__zz_execute_BranchPlugin_missAlignedTarget_6;
  wire       [31:0]   _zz__zz_execute_BranchPlugin_missAlignedTarget_6_1;
  wire       [31:0]   _zz__zz_execute_BranchPlugin_missAlignedTarget_6_2;
  wire       [19:0]   _zz__zz_execute_BranchPlugin_branch_src2_2;
  wire       [11:0]   _zz__zz_execute_BranchPlugin_branch_src2_4;
  wire                _zz_execute_BranchPlugin_branch_src2_6;
  wire                _zz_execute_BranchPlugin_branch_src2_7;
  wire                _zz_execute_BranchPlugin_branch_src2_8;
  wire       [2:0]    _zz_execute_BranchPlugin_branch_src2_9;
  wire       [1:0]    _zz__zz_CsrPlugin_exceptionPortCtrl_exceptionContext_code_1;
  wire       [1:0]    _zz__zz_CsrPlugin_exceptionPortCtrl_exceptionContext_code_1_1;
  wire                _zz_when;
  wire       [65:0]   _zz_writeBack_MulPlugin_result;
  wire       [65:0]   _zz_writeBack_MulPlugin_result_1;
  wire       [31:0]   _zz__zz_decode_RS2_2;
  wire       [31:0]   _zz__zz_decode_RS2_2_1;
  wire       [5:0]    _zz_memory_DivPlugin_div_counter_valueNext;
  wire       [0:0]    _zz_memory_DivPlugin_div_counter_valueNext_1;
  wire       [32:0]   _zz_memory_DivPlugin_div_stage_0_remainderMinusDenominator;
  wire       [31:0]   _zz_memory_DivPlugin_div_stage_0_outRemainder;
  wire       [31:0]   _zz_memory_DivPlugin_div_stage_0_outRemainder_1;
  wire       [32:0]   _zz_memory_DivPlugin_div_stage_0_outNumerator;
  wire       [32:0]   _zz_memory_DivPlugin_div_result_1;
  wire       [32:0]   _zz_memory_DivPlugin_div_result_2;
  wire       [32:0]   _zz_memory_DivPlugin_div_result_3;
  wire       [32:0]   _zz_memory_DivPlugin_div_result_4;
  wire       [0:0]    _zz_memory_DivPlugin_div_result_5;
  wire       [32:0]   _zz_memory_DivPlugin_rs1_2;
  wire       [0:0]    _zz_memory_DivPlugin_rs1_3;
  wire       [31:0]   _zz_memory_DivPlugin_rs2_1;
  wire       [0:0]    _zz_memory_DivPlugin_rs2_2;
  wire       [31:0]   _zz_PmpPlugin_pmpaddr_port;
  reg        [7:0]    _zz_when_PmpPlugin_l209;
  wire       [3:0]    _zz_when_PmpPlugin_l209_1;
  reg        [7:0]    _zz_when_PmpPlugin_l209_1_1;
  wire       [3:0]    _zz_when_PmpPlugin_l209_1_2;
  reg        [7:0]    _zz_when_PmpPlugin_l209_2;
  wire       [3:0]    _zz_when_PmpPlugin_l209_2_1;
  reg        [7:0]    _zz_when_PmpPlugin_l209_3;
  wire       [3:0]    _zz_when_PmpPlugin_l209_3_1;
  reg        [7:0]    _zz_when_PmpPlugin_l216;
  wire       [31:0]   _zz_CsrPlugin_csrMapping_readDataInit_25;
  reg        [7:0]    _zz_CsrPlugin_csrMapping_readDataSignal;
  wire       [3:0]    _zz_CsrPlugin_csrMapping_readDataSignal_1;
  reg        [7:0]    _zz_CsrPlugin_csrMapping_readDataSignal_2;
  wire       [3:0]    _zz_CsrPlugin_csrMapping_readDataSignal_3;
  reg        [7:0]    _zz_CsrPlugin_csrMapping_readDataSignal_4;
  wire       [3:0]    _zz_CsrPlugin_csrMapping_readDataSignal_5;
  reg        [7:0]    _zz_CsrPlugin_csrMapping_readDataSignal_6;
  wire       [3:0]    _zz_CsrPlugin_csrMapping_readDataSignal_7;
  wire       [26:0]   _zz_iBusWishbone_ADR_1;
  reg                 _zz_1;
  wire       [51:0]   memory_MUL_LOW;
  wire       [33:0]   memory_MUL_HH;
  wire       [33:0]   execute_MUL_HH;
  wire       [33:0]   execute_MUL_HL;
  wire       [33:0]   execute_MUL_LH;
  wire       [31:0]   execute_MUL_LL;
  wire       [31:0]   execute_BRANCH_CALC;
  wire                execute_BRANCH_DO;
  wire       [31:0]   execute_SHIFT_RIGHT;
  wire       [31:0]   execute_REGFILE_WRITE_DATA;
  wire       [31:0]   memory_MEMORY_STORE_DATA_RF;
  wire       [31:0]   execute_MEMORY_STORE_DATA_RF;
  wire                decode_CSR_READ_OPCODE;
  wire                decode_CSR_WRITE_OPCODE;
  wire                decode_PREDICTION_HAD_BRANCHED2;
  wire                decode_SRC2_FORCE_ZERO;
  wire                decode_IS_RS2_SIGNED;
  wire                decode_IS_RS1_SIGNED;
  wire                decode_IS_DIV;
  wire                memory_IS_MUL;
  wire                execute_IS_MUL;
  wire                decode_IS_MUL;
  wire       [1:0]    _zz_memory_to_writeBack_ENV_CTRL;
  wire       [1:0]    _zz_memory_to_writeBack_ENV_CTRL_1;
  wire       [1:0]    _zz_execute_to_memory_ENV_CTRL;
  wire       [1:0]    _zz_execute_to_memory_ENV_CTRL_1;
  wire       [1:0]    decode_ENV_CTRL;
  wire       [1:0]    _zz_decode_ENV_CTRL;
  wire       [1:0]    _zz_decode_to_execute_ENV_CTRL;
  wire       [1:0]    _zz_decode_to_execute_ENV_CTRL_1;
  wire                decode_IS_CSR;
  wire       [1:0]    _zz_decode_to_execute_BRANCH_CTRL;
  wire       [1:0]    _zz_decode_to_execute_BRANCH_CTRL_1;
  wire       [1:0]    _zz_execute_to_memory_SHIFT_CTRL;
  wire       [1:0]    _zz_execute_to_memory_SHIFT_CTRL_1;
  wire       [1:0]    decode_SHIFT_CTRL;
  wire       [1:0]    _zz_decode_SHIFT_CTRL;
  wire       [1:0]    _zz_decode_to_execute_SHIFT_CTRL;
  wire       [1:0]    _zz_decode_to_execute_SHIFT_CTRL_1;
  wire       [1:0]    decode_ALU_BITWISE_CTRL;
  wire       [1:0]    _zz_decode_ALU_BITWISE_CTRL;
  wire       [1:0]    _zz_decode_to_execute_ALU_BITWISE_CTRL;
  wire       [1:0]    _zz_decode_to_execute_ALU_BITWISE_CTRL_1;
  wire                decode_SRC_LESS_UNSIGNED;
  wire                decode_MEMORY_MANAGMENT;
  wire                memory_MEMORY_WR;
  wire                decode_MEMORY_WR;
  wire                execute_BYPASSABLE_MEMORY_STAGE;
  wire                decode_BYPASSABLE_MEMORY_STAGE;
  wire                decode_BYPASSABLE_EXECUTE_STAGE;
  wire       [1:0]    decode_SRC2_CTRL;
  wire       [1:0]    _zz_decode_SRC2_CTRL;
  wire       [1:0]    _zz_decode_to_execute_SRC2_CTRL;
  wire       [1:0]    _zz_decode_to_execute_SRC2_CTRL_1;
  wire       [1:0]    decode_ALU_CTRL;
  wire       [1:0]    _zz_decode_ALU_CTRL;
  wire       [1:0]    _zz_decode_to_execute_ALU_CTRL;
  wire       [1:0]    _zz_decode_to_execute_ALU_CTRL_1;
  wire       [1:0]    decode_SRC1_CTRL;
  wire       [1:0]    _zz_decode_SRC1_CTRL;
  wire       [1:0]    _zz_decode_to_execute_SRC1_CTRL;
  wire       [1:0]    _zz_decode_to_execute_SRC1_CTRL_1;
  wire                decode_MEMORY_FORCE_CONSTISTENCY;
  wire       [31:0]   writeBack_FORMAL_PC_NEXT;
  wire       [31:0]   memory_FORMAL_PC_NEXT;
  wire       [31:0]   execute_FORMAL_PC_NEXT;
  wire       [31:0]   decode_FORMAL_PC_NEXT;
  wire       [31:0]   memory_PC;
  wire                execute_IS_RS1_SIGNED;
  wire                execute_IS_DIV;
  wire                execute_IS_RS2_SIGNED;
  wire                memory_IS_DIV;
  wire                writeBack_IS_MUL;
  wire       [33:0]   writeBack_MUL_HH;
  wire       [51:0]   writeBack_MUL_LOW;
  wire       [33:0]   memory_MUL_HL;
  wire       [33:0]   memory_MUL_LH;
  wire       [31:0]   memory_MUL_LL;
  wire                execute_CSR_READ_OPCODE;
  wire                execute_CSR_WRITE_OPCODE;
  wire                execute_IS_CSR;
  wire       [1:0]    memory_ENV_CTRL;
  wire       [1:0]    _zz_memory_ENV_CTRL;
  wire       [1:0]    execute_ENV_CTRL;
  wire       [1:0]    _zz_execute_ENV_CTRL;
  wire       [1:0]    writeBack_ENV_CTRL;
  wire       [1:0]    _zz_writeBack_ENV_CTRL;
  wire       [31:0]   memory_BRANCH_CALC;
  wire                memory_BRANCH_DO;
  wire       [31:0]   execute_PC;
  wire                execute_PREDICTION_HAD_BRANCHED2;
  wire                execute_BRANCH_COND_RESULT;
  wire       [1:0]    execute_BRANCH_CTRL;
  wire       [1:0]    _zz_execute_BRANCH_CTRL;
  wire                decode_RS2_USE;
  wire                decode_RS1_USE;
  reg        [31:0]   _zz_decode_RS2;
  wire                execute_REGFILE_WRITE_VALID;
  wire                execute_BYPASSABLE_EXECUTE_STAGE;
  wire                memory_REGFILE_WRITE_VALID;
  wire       [31:0]   memory_INSTRUCTION;
  wire                memory_BYPASSABLE_MEMORY_STAGE;
  wire                writeBack_REGFILE_WRITE_VALID;
  reg        [31:0]   decode_RS2;
  reg        [31:0]   decode_RS1;
  wire       [31:0]   memory_SHIFT_RIGHT;
  reg        [31:0]   _zz_decode_RS2_1;
  wire       [1:0]    memory_SHIFT_CTRL;
  wire       [1:0]    _zz_memory_SHIFT_CTRL;
  wire       [1:0]    execute_SHIFT_CTRL;
  wire       [1:0]    _zz_execute_SHIFT_CTRL;
  wire                execute_SRC_LESS_UNSIGNED;
  wire                execute_SRC2_FORCE_ZERO;
  wire                execute_SRC_USE_SUB_LESS;
  wire       [31:0]   _zz_execute_SRC2;
  wire       [1:0]    execute_SRC2_CTRL;
  wire       [1:0]    _zz_execute_SRC2_CTRL;
  wire       [1:0]    execute_SRC1_CTRL;
  wire       [1:0]    _zz_execute_SRC1_CTRL;
  wire                decode_SRC_USE_SUB_LESS;
  wire                decode_SRC_ADD_ZERO;
  wire       [31:0]   execute_SRC_ADD_SUB;
  wire                execute_SRC_LESS;
  wire       [1:0]    execute_ALU_CTRL;
  wire       [1:0]    _zz_execute_ALU_CTRL;
  wire       [31:0]   execute_SRC2;
  wire       [31:0]   execute_SRC1;
  wire       [1:0]    execute_ALU_BITWISE_CTRL;
  wire       [1:0]    _zz_execute_ALU_BITWISE_CTRL;
  wire       [31:0]   _zz_lastStageRegFileWrite_payload_address;
  wire                _zz_lastStageRegFileWrite_valid;
  reg                 _zz_2;
  wire       [31:0]   decode_INSTRUCTION_ANTICIPATED;
  reg                 decode_REGFILE_WRITE_VALID;
  wire                decode_LEGAL_INSTRUCTION;
  wire       [1:0]    _zz_decode_ENV_CTRL_1;
  wire       [1:0]    _zz_decode_BRANCH_CTRL;
  wire       [1:0]    _zz_decode_SHIFT_CTRL_1;
  wire       [1:0]    _zz_decode_ALU_BITWISE_CTRL_1;
  wire       [1:0]    _zz_decode_SRC2_CTRL_1;
  wire       [1:0]    _zz_decode_ALU_CTRL_1;
  wire       [1:0]    _zz_decode_SRC1_CTRL_1;
  reg        [31:0]   _zz_decode_RS2_2;
  wire                writeBack_MEMORY_WR;
  wire       [31:0]   writeBack_MEMORY_STORE_DATA_RF;
  wire       [31:0]   writeBack_REGFILE_WRITE_DATA;
  wire                writeBack_MEMORY_ENABLE;
  wire       [31:0]   memory_REGFILE_WRITE_DATA;
  wire                memory_MEMORY_ENABLE;
  wire                execute_MEMORY_FORCE_CONSTISTENCY;
  (* keep , syn_keep *) wire       [31:0]   execute_RS1 /* synthesis syn_keep = 1 */ ;
  wire                execute_MEMORY_MANAGMENT;
  (* keep , syn_keep *) wire       [31:0]   execute_RS2 /* synthesis syn_keep = 1 */ ;
  wire                execute_MEMORY_WR;
  wire       [31:0]   execute_SRC_ADD;
  wire                execute_MEMORY_ENABLE;
  wire       [31:0]   execute_INSTRUCTION;
  wire                decode_MEMORY_ENABLE;
  wire                decode_FLUSH_ALL;
  reg                 IBusCachedPlugin_rsp_issueDetected_4;
  reg                 IBusCachedPlugin_rsp_issueDetected_3;
  reg                 IBusCachedPlugin_rsp_issueDetected_2;
  reg                 IBusCachedPlugin_rsp_issueDetected_1;
  wire       [1:0]    decode_BRANCH_CTRL;
  wire       [1:0]    _zz_decode_BRANCH_CTRL_1;
  wire       [31:0]   decode_INSTRUCTION;
  reg        [31:0]   _zz_memory_to_writeBack_FORMAL_PC_NEXT;
  reg        [31:0]   _zz_decode_to_execute_FORMAL_PC_NEXT;
  wire       [31:0]   decode_PC;
  wire       [31:0]   writeBack_PC;
  wire       [31:0]   writeBack_INSTRUCTION;
  reg                 decode_arbitration_haltItself;
  reg                 decode_arbitration_haltByOther;
  reg                 decode_arbitration_removeIt;
  wire                decode_arbitration_flushIt;
  reg                 decode_arbitration_flushNext;
  reg                 decode_arbitration_isValid;
  wire                decode_arbitration_isStuck;
  wire                decode_arbitration_isStuckByOthers;
  wire                decode_arbitration_isFlushed;
  wire                decode_arbitration_isMoving;
  wire                decode_arbitration_isFiring;
  reg                 execute_arbitration_haltItself;
  reg                 execute_arbitration_haltByOther;
  reg                 execute_arbitration_removeIt;
  wire                execute_arbitration_flushIt;
  reg                 execute_arbitration_flushNext;
  reg                 execute_arbitration_isValid;
  wire                execute_arbitration_isStuck;
  wire                execute_arbitration_isStuckByOthers;
  wire                execute_arbitration_isFlushed;
  wire                execute_arbitration_isMoving;
  wire                execute_arbitration_isFiring;
  reg                 memory_arbitration_haltItself;
  wire                memory_arbitration_haltByOther;
  reg                 memory_arbitration_removeIt;
  wire                memory_arbitration_flushIt;
  reg                 memory_arbitration_flushNext;
  reg                 memory_arbitration_isValid;
  wire                memory_arbitration_isStuck;
  wire                memory_arbitration_isStuckByOthers;
  wire                memory_arbitration_isFlushed;
  wire                memory_arbitration_isMoving;
  wire                memory_arbitration_isFiring;
  reg                 writeBack_arbitration_haltItself;
  wire                writeBack_arbitration_haltByOther;
  reg                 writeBack_arbitration_removeIt;
  reg                 writeBack_arbitration_flushIt;
  reg                 writeBack_arbitration_flushNext;
  reg                 writeBack_arbitration_isValid;
  wire                writeBack_arbitration_isStuck;
  wire                writeBack_arbitration_isStuckByOthers;
  wire                writeBack_arbitration_isFlushed;
  wire                writeBack_arbitration_isMoving;
  wire                writeBack_arbitration_isFiring;
  wire       [31:0]   lastStageInstruction /* verilator public */ ;
  wire       [31:0]   lastStagePc /* verilator public */ ;
  wire                lastStageIsValid /* verilator public */ ;
  wire                lastStageIsFiring /* verilator public */ ;
  reg                 IBusCachedPlugin_fetcherHalt;
  wire                IBusCachedPlugin_forceNoDecodeCond;
  reg                 IBusCachedPlugin_incomingInstruction;
  wire                IBusCachedPlugin_predictionJumpInterface_valid;
  (* keep , syn_keep *) wire       [31:0]   IBusCachedPlugin_predictionJumpInterface_payload /* synthesis syn_keep = 1 */ ;
  reg                 IBusCachedPlugin_decodePrediction_cmd_hadBranch;
  wire                IBusCachedPlugin_decodePrediction_rsp_wasWrong;
  wire                IBusCachedPlugin_pcValids_0;
  wire                IBusCachedPlugin_pcValids_1;
  wire                IBusCachedPlugin_pcValids_2;
  wire                IBusCachedPlugin_pcValids_3;
  reg                 IBusCachedPlugin_decodeExceptionPort_valid;
  reg        [3:0]    IBusCachedPlugin_decodeExceptionPort_payload_code;
  wire       [31:0]   IBusCachedPlugin_decodeExceptionPort_payload_badAddr;
  wire                IBusCachedPlugin_mmuBus_cmd_0_isValid;
  wire                IBusCachedPlugin_mmuBus_cmd_0_isStuck;
  wire       [31:0]   IBusCachedPlugin_mmuBus_cmd_0_virtualAddress;
  wire                IBusCachedPlugin_mmuBus_cmd_0_bypassTranslation;
  wire       [31:0]   IBusCachedPlugin_mmuBus_rsp_physicalAddress;
  wire                IBusCachedPlugin_mmuBus_rsp_isIoAccess;
  wire                IBusCachedPlugin_mmuBus_rsp_isPaging;
  wire                IBusCachedPlugin_mmuBus_rsp_allowRead;
  wire                IBusCachedPlugin_mmuBus_rsp_allowWrite;
  reg                 IBusCachedPlugin_mmuBus_rsp_allowExecute;
  wire                IBusCachedPlugin_mmuBus_rsp_exception;
  wire                IBusCachedPlugin_mmuBus_rsp_refilling;
  wire                IBusCachedPlugin_mmuBus_rsp_bypassTranslation;
  wire                IBusCachedPlugin_mmuBus_end;
  wire                IBusCachedPlugin_mmuBus_busy;
  wire                dBus_cmd_valid;
  wire                dBus_cmd_ready;
  wire                dBus_cmd_payload_wr;
  wire                dBus_cmd_payload_uncached;
  wire       [31:0]   dBus_cmd_payload_address;
  wire       [31:0]   dBus_cmd_payload_data;
  wire       [3:0]    dBus_cmd_payload_mask;
  wire       [2:0]    dBus_cmd_payload_size;
  wire                dBus_cmd_payload_last;
  wire                dBus_rsp_valid;
  wire                dBus_rsp_payload_last;
  wire       [31:0]   dBus_rsp_payload_data;
  wire                dBus_rsp_payload_error;
  wire                DBusCachedPlugin_mmuBus_cmd_0_isValid;
  wire                DBusCachedPlugin_mmuBus_cmd_0_isStuck;
  wire       [31:0]   DBusCachedPlugin_mmuBus_cmd_0_virtualAddress;
  wire                DBusCachedPlugin_mmuBus_cmd_0_bypassTranslation;
  wire       [31:0]   DBusCachedPlugin_mmuBus_rsp_physicalAddress;
  wire                DBusCachedPlugin_mmuBus_rsp_isIoAccess;
  wire                DBusCachedPlugin_mmuBus_rsp_isPaging;
  reg                 DBusCachedPlugin_mmuBus_rsp_allowRead;
  reg                 DBusCachedPlugin_mmuBus_rsp_allowWrite;
  wire                DBusCachedPlugin_mmuBus_rsp_allowExecute;
  wire                DBusCachedPlugin_mmuBus_rsp_exception;
  wire                DBusCachedPlugin_mmuBus_rsp_refilling;
  wire                DBusCachedPlugin_mmuBus_rsp_bypassTranslation;
  wire                DBusCachedPlugin_mmuBus_end;
  wire                DBusCachedPlugin_mmuBus_busy;
  reg                 DBusCachedPlugin_redoBranch_valid;
  wire       [31:0]   DBusCachedPlugin_redoBranch_payload;
  reg                 DBusCachedPlugin_exceptionBus_valid;
  reg        [3:0]    DBusCachedPlugin_exceptionBus_payload_code;
  wire       [31:0]   DBusCachedPlugin_exceptionBus_payload_badAddr;
  wire                decodeExceptionPort_valid;
  wire       [3:0]    decodeExceptionPort_payload_code;
  wire       [31:0]   decodeExceptionPort_payload_badAddr;
  wire                BranchPlugin_jumpInterface_valid;
  wire       [31:0]   BranchPlugin_jumpInterface_payload;
  wire                BranchPlugin_branchExceptionPort_valid;
  wire       [3:0]    BranchPlugin_branchExceptionPort_payload_code;
  wire       [31:0]   BranchPlugin_branchExceptionPort_payload_badAddr;
  wire                BranchPlugin_inDebugNoFetchFlag;
  reg        [31:0]   CsrPlugin_csrMapping_readDataSignal;
  wire       [31:0]   CsrPlugin_csrMapping_readDataInit;
  wire       [31:0]   CsrPlugin_csrMapping_writeDataSignal;
  reg                 CsrPlugin_csrMapping_allowCsrSignal;
  wire                CsrPlugin_csrMapping_hazardFree;
  reg                 CsrPlugin_inWfi /* verilator public */ ;
  wire                CsrPlugin_thirdPartyWake;
  reg                 CsrPlugin_jumpInterface_valid;
  reg        [31:0]   CsrPlugin_jumpInterface_payload;
  wire                CsrPlugin_exceptionPendings_0;
  wire                CsrPlugin_exceptionPendings_1;
  wire                CsrPlugin_exceptionPendings_2;
  wire                CsrPlugin_exceptionPendings_3;
  wire                externalInterrupt;
  wire                contextSwitching;
  reg        [1:0]    CsrPlugin_privilege;
  wire                CsrPlugin_forceMachineWire;
  reg                 CsrPlugin_selfException_valid;
  reg        [3:0]    CsrPlugin_selfException_payload_code;
  wire       [31:0]   CsrPlugin_selfException_payload_badAddr;
  wire                CsrPlugin_allowInterrupts;
  wire                CsrPlugin_allowException;
  wire                CsrPlugin_allowEbreakException;
  wire                IBusCachedPlugin_externalFlush;
  wire                IBusCachedPlugin_jump_pcLoad_valid;
  wire       [31:0]   IBusCachedPlugin_jump_pcLoad_payload;
  wire       [3:0]    _zz_IBusCachedPlugin_jump_pcLoad_payload;
  wire       [3:0]    _zz_IBusCachedPlugin_jump_pcLoad_payload_1;
  wire                _zz_IBusCachedPlugin_jump_pcLoad_payload_2;
  wire                _zz_IBusCachedPlugin_jump_pcLoad_payload_3;
  wire                _zz_IBusCachedPlugin_jump_pcLoad_payload_4;
  wire                IBusCachedPlugin_fetchPc_output_valid;
  wire                IBusCachedPlugin_fetchPc_output_ready;
  wire       [31:0]   IBusCachedPlugin_fetchPc_output_payload;
  reg        [31:0]   IBusCachedPlugin_fetchPc_pcReg /* verilator public */ ;
  reg                 IBusCachedPlugin_fetchPc_correction;
  reg                 IBusCachedPlugin_fetchPc_correctionReg;
  wire                IBusCachedPlugin_fetchPc_output_fire;
  wire                IBusCachedPlugin_fetchPc_corrected;
  reg                 IBusCachedPlugin_fetchPc_pcRegPropagate;
  reg                 IBusCachedPlugin_fetchPc_booted;
  reg                 IBusCachedPlugin_fetchPc_inc;
  wire                when_Fetcher_l134;
  wire                IBusCachedPlugin_fetchPc_output_fire_1;
  wire                when_Fetcher_l134_1;
  reg        [31:0]   IBusCachedPlugin_fetchPc_pc;
  wire                IBusCachedPlugin_fetchPc_redo_valid;
  wire       [31:0]   IBusCachedPlugin_fetchPc_redo_payload;
  reg                 IBusCachedPlugin_fetchPc_flushed;
  wire                when_Fetcher_l161;
  reg                 IBusCachedPlugin_iBusRsp_redoFetch;
  wire                IBusCachedPlugin_iBusRsp_stages_0_input_valid;
  wire                IBusCachedPlugin_iBusRsp_stages_0_input_ready;
  wire       [31:0]   IBusCachedPlugin_iBusRsp_stages_0_input_payload;
  wire                IBusCachedPlugin_iBusRsp_stages_0_output_valid;
  wire                IBusCachedPlugin_iBusRsp_stages_0_output_ready;
  wire       [31:0]   IBusCachedPlugin_iBusRsp_stages_0_output_payload;
  reg                 IBusCachedPlugin_iBusRsp_stages_0_halt;
  wire                IBusCachedPlugin_iBusRsp_stages_1_input_valid;
  wire                IBusCachedPlugin_iBusRsp_stages_1_input_ready;
  wire       [31:0]   IBusCachedPlugin_iBusRsp_stages_1_input_payload;
  wire                IBusCachedPlugin_iBusRsp_stages_1_output_valid;
  wire                IBusCachedPlugin_iBusRsp_stages_1_output_ready;
  wire       [31:0]   IBusCachedPlugin_iBusRsp_stages_1_output_payload;
  reg                 IBusCachedPlugin_iBusRsp_stages_1_halt;
  wire                IBusCachedPlugin_iBusRsp_stages_2_input_valid;
  wire                IBusCachedPlugin_iBusRsp_stages_2_input_ready;
  wire       [31:0]   IBusCachedPlugin_iBusRsp_stages_2_input_payload;
  wire                IBusCachedPlugin_iBusRsp_stages_2_output_valid;
  wire                IBusCachedPlugin_iBusRsp_stages_2_output_ready;
  wire       [31:0]   IBusCachedPlugin_iBusRsp_stages_2_output_payload;
  reg                 IBusCachedPlugin_iBusRsp_stages_2_halt;
  wire                _zz_IBusCachedPlugin_iBusRsp_stages_0_input_ready;
  wire                _zz_IBusCachedPlugin_iBusRsp_stages_1_input_ready;
  wire                _zz_IBusCachedPlugin_iBusRsp_stages_2_input_ready;
  wire                IBusCachedPlugin_iBusRsp_flush;
  wire                _zz_IBusCachedPlugin_iBusRsp_stages_0_output_ready;
  wire                _zz_IBusCachedPlugin_iBusRsp_stages_0_output_ready_1;
  reg                 _zz_IBusCachedPlugin_iBusRsp_stages_0_output_ready_2;
  wire                IBusCachedPlugin_iBusRsp_stages_1_output_m2sPipe_valid;
  wire                IBusCachedPlugin_iBusRsp_stages_1_output_m2sPipe_ready;
  wire       [31:0]   IBusCachedPlugin_iBusRsp_stages_1_output_m2sPipe_payload;
  reg                 _zz_IBusCachedPlugin_iBusRsp_stages_1_output_m2sPipe_valid;
  reg        [31:0]   _zz_IBusCachedPlugin_iBusRsp_stages_1_output_m2sPipe_payload;
  reg                 IBusCachedPlugin_iBusRsp_readyForError;
  wire                IBusCachedPlugin_iBusRsp_output_valid;
  wire                IBusCachedPlugin_iBusRsp_output_ready;
  wire       [31:0]   IBusCachedPlugin_iBusRsp_output_payload_pc;
  wire                IBusCachedPlugin_iBusRsp_output_payload_rsp_error;
  wire       [31:0]   IBusCachedPlugin_iBusRsp_output_payload_rsp_inst;
  wire                IBusCachedPlugin_iBusRsp_output_payload_isRvc;
  wire                when_Fetcher_l243;
  wire                when_Fetcher_l323;
  reg                 IBusCachedPlugin_injector_nextPcCalc_valids_0;
  wire                when_Fetcher_l332;
  reg                 IBusCachedPlugin_injector_nextPcCalc_valids_1;
  wire                when_Fetcher_l332_1;
  reg                 IBusCachedPlugin_injector_nextPcCalc_valids_2;
  wire                when_Fetcher_l332_2;
  reg                 IBusCachedPlugin_injector_nextPcCalc_valids_3;
  wire                when_Fetcher_l332_3;
  reg                 IBusCachedPlugin_injector_nextPcCalc_valids_4;
  wire                when_Fetcher_l332_4;
  wire                _zz_IBusCachedPlugin_decodePrediction_cmd_hadBranch;
  reg        [18:0]   _zz_IBusCachedPlugin_decodePrediction_cmd_hadBranch_1;
  wire                _zz_3;
  reg        [10:0]   _zz_4;
  wire                _zz_5;
  reg        [18:0]   _zz_6;
  reg                 _zz_7;
  wire                _zz_IBusCachedPlugin_predictionJumpInterface_payload;
  reg        [10:0]   _zz_IBusCachedPlugin_predictionJumpInterface_payload_1;
  wire                _zz_IBusCachedPlugin_predictionJumpInterface_payload_2;
  reg        [18:0]   _zz_IBusCachedPlugin_predictionJumpInterface_payload_3;
  wire                iBus_cmd_valid;
  wire                iBus_cmd_ready;
  reg        [31:0]   iBus_cmd_payload_address;
  wire       [2:0]    iBus_cmd_payload_size;
  wire                iBus_rsp_valid;
  wire       [31:0]   iBus_rsp_payload_data;
  wire                iBus_rsp_payload_error;
  reg        [31:0]   IBusCachedPlugin_rspCounter;
  wire                IBusCachedPlugin_s0_tightlyCoupledHit;
  reg                 IBusCachedPlugin_s1_tightlyCoupledHit;
  reg                 IBusCachedPlugin_s2_tightlyCoupledHit;
  wire                IBusCachedPlugin_rsp_iBusRspOutputHalt;
  wire                IBusCachedPlugin_rsp_issueDetected;
  reg                 IBusCachedPlugin_rsp_redoFetch;
  wire                when_IBusCachedPlugin_l239;
  wire                when_IBusCachedPlugin_l244;
  wire                when_IBusCachedPlugin_l250;
  wire                when_IBusCachedPlugin_l256;
  wire                when_IBusCachedPlugin_l267;
  wire                dataCache_1_io_mem_cmd_s2mPipe_valid;
  reg                 dataCache_1_io_mem_cmd_s2mPipe_ready;
  wire                dataCache_1_io_mem_cmd_s2mPipe_payload_wr;
  wire                dataCache_1_io_mem_cmd_s2mPipe_payload_uncached;
  wire       [31:0]   dataCache_1_io_mem_cmd_s2mPipe_payload_address;
  wire       [31:0]   dataCache_1_io_mem_cmd_s2mPipe_payload_data;
  wire       [3:0]    dataCache_1_io_mem_cmd_s2mPipe_payload_mask;
  wire       [2:0]    dataCache_1_io_mem_cmd_s2mPipe_payload_size;
  wire                dataCache_1_io_mem_cmd_s2mPipe_payload_last;
  reg                 dataCache_1_io_mem_cmd_rValid;
  reg                 dataCache_1_io_mem_cmd_rData_wr;
  reg                 dataCache_1_io_mem_cmd_rData_uncached;
  reg        [31:0]   dataCache_1_io_mem_cmd_rData_address;
  reg        [31:0]   dataCache_1_io_mem_cmd_rData_data;
  reg        [3:0]    dataCache_1_io_mem_cmd_rData_mask;
  reg        [2:0]    dataCache_1_io_mem_cmd_rData_size;
  reg                 dataCache_1_io_mem_cmd_rData_last;
  wire                dataCache_1_io_mem_cmd_s2mPipe_m2sPipe_valid;
  wire                dataCache_1_io_mem_cmd_s2mPipe_m2sPipe_ready;
  wire                dataCache_1_io_mem_cmd_s2mPipe_m2sPipe_payload_wr;
  wire                dataCache_1_io_mem_cmd_s2mPipe_m2sPipe_payload_uncached;
  wire       [31:0]   dataCache_1_io_mem_cmd_s2mPipe_m2sPipe_payload_address;
  wire       [31:0]   dataCache_1_io_mem_cmd_s2mPipe_m2sPipe_payload_data;
  wire       [3:0]    dataCache_1_io_mem_cmd_s2mPipe_m2sPipe_payload_mask;
  wire       [2:0]    dataCache_1_io_mem_cmd_s2mPipe_m2sPipe_payload_size;
  wire                dataCache_1_io_mem_cmd_s2mPipe_m2sPipe_payload_last;
  reg                 dataCache_1_io_mem_cmd_s2mPipe_rValid;
  reg                 dataCache_1_io_mem_cmd_s2mPipe_rData_wr;
  reg                 dataCache_1_io_mem_cmd_s2mPipe_rData_uncached;
  reg        [31:0]   dataCache_1_io_mem_cmd_s2mPipe_rData_address;
  reg        [31:0]   dataCache_1_io_mem_cmd_s2mPipe_rData_data;
  reg        [3:0]    dataCache_1_io_mem_cmd_s2mPipe_rData_mask;
  reg        [2:0]    dataCache_1_io_mem_cmd_s2mPipe_rData_size;
  reg                 dataCache_1_io_mem_cmd_s2mPipe_rData_last;
  wire                when_Stream_l368;
  reg        [31:0]   DBusCachedPlugin_rspCounter;
  wire                when_DBusCachedPlugin_l308;
  wire       [1:0]    execute_DBusCachedPlugin_size;
  reg        [31:0]   _zz_execute_MEMORY_STORE_DATA_RF;
  wire                dataCache_1_io_cpu_flush_isStall;
  wire                when_DBusCachedPlugin_l350;
  wire                when_DBusCachedPlugin_l366;
  wire                when_DBusCachedPlugin_l393;
  wire                when_DBusCachedPlugin_l446;
  wire                when_DBusCachedPlugin_l466;
  wire       [7:0]    writeBack_DBusCachedPlugin_rspSplits_0;
  wire       [7:0]    writeBack_DBusCachedPlugin_rspSplits_1;
  wire       [7:0]    writeBack_DBusCachedPlugin_rspSplits_2;
  wire       [7:0]    writeBack_DBusCachedPlugin_rspSplits_3;
  reg        [31:0]   writeBack_DBusCachedPlugin_rspShifted;
  wire       [31:0]   writeBack_DBusCachedPlugin_rspRf;
  wire       [1:0]    switch_Misc_l210;
  wire                _zz_writeBack_DBusCachedPlugin_rspFormated;
  reg        [31:0]   _zz_writeBack_DBusCachedPlugin_rspFormated_1;
  wire                _zz_writeBack_DBusCachedPlugin_rspFormated_2;
  reg        [31:0]   _zz_writeBack_DBusCachedPlugin_rspFormated_3;
  reg        [31:0]   writeBack_DBusCachedPlugin_rspFormated;
  wire                when_DBusCachedPlugin_l492;
  reg        [7:0]    PmpPlugin_pmpcfg_0;
  reg        [7:0]    PmpPlugin_pmpcfg_1;
  reg        [7:0]    PmpPlugin_pmpcfg_2;
  reg        [7:0]    PmpPlugin_pmpcfg_3;
  reg        [7:0]    PmpPlugin_pmpcfg_4;
  reg        [7:0]    PmpPlugin_pmpcfg_5;
  reg        [7:0]    PmpPlugin_pmpcfg_6;
  reg        [7:0]    PmpPlugin_pmpcfg_7;
  reg        [7:0]    PmpPlugin_pmpcfg_8;
  reg        [7:0]    PmpPlugin_pmpcfg_9;
  reg        [7:0]    PmpPlugin_pmpcfg_10;
  reg        [7:0]    PmpPlugin_pmpcfg_11;
  reg        [7:0]    PmpPlugin_pmpcfg_12;
  reg        [7:0]    PmpPlugin_pmpcfg_13;
  reg        [7:0]    PmpPlugin_pmpcfg_14;
  reg        [7:0]    PmpPlugin_pmpcfg_15;
  reg        [24:0]   PmpPlugin_base_0;
  reg        [24:0]   PmpPlugin_base_1;
  reg        [24:0]   PmpPlugin_base_2;
  reg        [24:0]   PmpPlugin_base_3;
  reg        [24:0]   PmpPlugin_base_4;
  reg        [24:0]   PmpPlugin_base_5;
  reg        [24:0]   PmpPlugin_base_6;
  reg        [24:0]   PmpPlugin_base_7;
  reg        [24:0]   PmpPlugin_base_8;
  reg        [24:0]   PmpPlugin_base_9;
  reg        [24:0]   PmpPlugin_base_10;
  reg        [24:0]   PmpPlugin_base_11;
  reg        [24:0]   PmpPlugin_base_12;
  reg        [24:0]   PmpPlugin_base_13;
  reg        [24:0]   PmpPlugin_base_14;
  reg        [24:0]   PmpPlugin_base_15;
  reg        [24:0]   PmpPlugin_mask_0;
  reg        [24:0]   PmpPlugin_mask_1;
  reg        [24:0]   PmpPlugin_mask_2;
  reg        [24:0]   PmpPlugin_mask_3;
  reg        [24:0]   PmpPlugin_mask_4;
  reg        [24:0]   PmpPlugin_mask_5;
  reg        [24:0]   PmpPlugin_mask_6;
  reg        [24:0]   PmpPlugin_mask_7;
  reg        [24:0]   PmpPlugin_mask_8;
  reg        [24:0]   PmpPlugin_mask_9;
  reg        [24:0]   PmpPlugin_mask_10;
  reg        [24:0]   PmpPlugin_mask_11;
  reg        [24:0]   PmpPlugin_mask_12;
  reg        [24:0]   PmpPlugin_mask_13;
  reg        [24:0]   PmpPlugin_mask_14;
  reg        [24:0]   PmpPlugin_mask_15;
  reg                 execute_PmpPlugin_fsmPending;
  wire                when_PmpPlugin_l138;
  reg                 execute_PmpPlugin_fsmComplete;
  wire       [11:0]   execute_PmpPlugin_csrAddress;
  wire       [3:0]    execute_PmpPlugin_pmpNcfg;
  wire       [1:0]    execute_PmpPlugin_pmpcfgN;
  wire                execute_PmpPlugin_pmpcfgCsr;
  wire                execute_PmpPlugin_pmpaddrCsr;
  reg        [3:0]    execute_PmpPlugin_pmpNcfg_;
  reg        [1:0]    execute_PmpPlugin_pmpcfgN_;
  reg                 execute_PmpPlugin_pmpcfgCsr_;
  reg                 execute_PmpPlugin_pmpaddrCsr_;
  reg        [31:0]   execute_PmpPlugin_writeData_;
  wire                execute_PmpPlugin_fsm_wantExit;
  reg                 execute_PmpPlugin_fsm_wantStart;
  wire                execute_PmpPlugin_fsm_wantKill;
  reg                 execute_PmpPlugin_fsm_fsmEnable;
  reg        [3:0]    execute_PmpPlugin_fsm_fsmCounter;
  wire                when_PmpPlugin_l246;
  wire       [15:0]   _zz_8;
  wire       [15:0]   _zz_9;
  wire       [24:0]   _zz_PmpPlugin_dGuard_hits_0;
  wire                PmpPlugin_dGuard_hits_0;
  wire                PmpPlugin_dGuard_hits_1;
  wire                PmpPlugin_dGuard_hits_2;
  wire                PmpPlugin_dGuard_hits_3;
  wire                PmpPlugin_dGuard_hits_4;
  wire                PmpPlugin_dGuard_hits_5;
  wire                PmpPlugin_dGuard_hits_6;
  wire                PmpPlugin_dGuard_hits_7;
  wire                PmpPlugin_dGuard_hits_8;
  wire                PmpPlugin_dGuard_hits_9;
  wire                PmpPlugin_dGuard_hits_10;
  wire                PmpPlugin_dGuard_hits_11;
  wire                PmpPlugin_dGuard_hits_12;
  wire                PmpPlugin_dGuard_hits_13;
  wire                PmpPlugin_dGuard_hits_14;
  wire                PmpPlugin_dGuard_hits_15;
  wire                when_PmpPlugin_l277;
  wire       [15:0]   _zz_DBusCachedPlugin_mmuBus_rsp_allowRead;
  wire       [15:0]   _zz_DBusCachedPlugin_mmuBus_rsp_allowRead_1;
  wire                _zz_DBusCachedPlugin_mmuBus_rsp_allowRead_2;
  wire                _zz_DBusCachedPlugin_mmuBus_rsp_allowRead_3;
  wire                _zz_DBusCachedPlugin_mmuBus_rsp_allowRead_4;
  wire                _zz_DBusCachedPlugin_mmuBus_rsp_allowRead_5;
  wire                _zz_DBusCachedPlugin_mmuBus_rsp_allowRead_6;
  wire                _zz_DBusCachedPlugin_mmuBus_rsp_allowRead_7;
  wire                _zz_DBusCachedPlugin_mmuBus_rsp_allowRead_8;
  wire                _zz_DBusCachedPlugin_mmuBus_rsp_allowRead_9;
  wire                _zz_DBusCachedPlugin_mmuBus_rsp_allowRead_10;
  wire                _zz_DBusCachedPlugin_mmuBus_rsp_allowRead_11;
  wire                _zz_DBusCachedPlugin_mmuBus_rsp_allowRead_12;
  wire                _zz_DBusCachedPlugin_mmuBus_rsp_allowRead_13;
  wire                _zz_DBusCachedPlugin_mmuBus_rsp_allowRead_14;
  wire                _zz_DBusCachedPlugin_mmuBus_rsp_allowRead_15;
  wire                _zz_DBusCachedPlugin_mmuBus_rsp_allowRead_16;
  wire       [15:0]   _zz_DBusCachedPlugin_mmuBus_rsp_allowWrite;
  wire       [15:0]   _zz_DBusCachedPlugin_mmuBus_rsp_allowWrite_1;
  wire                _zz_DBusCachedPlugin_mmuBus_rsp_allowWrite_2;
  wire                _zz_DBusCachedPlugin_mmuBus_rsp_allowWrite_3;
  wire                _zz_DBusCachedPlugin_mmuBus_rsp_allowWrite_4;
  wire                _zz_DBusCachedPlugin_mmuBus_rsp_allowWrite_5;
  wire                _zz_DBusCachedPlugin_mmuBus_rsp_allowWrite_6;
  wire                _zz_DBusCachedPlugin_mmuBus_rsp_allowWrite_7;
  wire                _zz_DBusCachedPlugin_mmuBus_rsp_allowWrite_8;
  wire                _zz_DBusCachedPlugin_mmuBus_rsp_allowWrite_9;
  wire                _zz_DBusCachedPlugin_mmuBus_rsp_allowWrite_10;
  wire                _zz_DBusCachedPlugin_mmuBus_rsp_allowWrite_11;
  wire                _zz_DBusCachedPlugin_mmuBus_rsp_allowWrite_12;
  wire                _zz_DBusCachedPlugin_mmuBus_rsp_allowWrite_13;
  wire                _zz_DBusCachedPlugin_mmuBus_rsp_allowWrite_14;
  wire                _zz_DBusCachedPlugin_mmuBus_rsp_allowWrite_15;
  wire                _zz_DBusCachedPlugin_mmuBus_rsp_allowWrite_16;
  wire       [24:0]   _zz_PmpPlugin_iGuard_hits_0;
  wire                PmpPlugin_iGuard_hits_0;
  wire                PmpPlugin_iGuard_hits_1;
  wire                PmpPlugin_iGuard_hits_2;
  wire                PmpPlugin_iGuard_hits_3;
  wire                PmpPlugin_iGuard_hits_4;
  wire                PmpPlugin_iGuard_hits_5;
  wire                PmpPlugin_iGuard_hits_6;
  wire                PmpPlugin_iGuard_hits_7;
  wire                PmpPlugin_iGuard_hits_8;
  wire                PmpPlugin_iGuard_hits_9;
  wire                PmpPlugin_iGuard_hits_10;
  wire                PmpPlugin_iGuard_hits_11;
  wire                PmpPlugin_iGuard_hits_12;
  wire                PmpPlugin_iGuard_hits_13;
  wire                PmpPlugin_iGuard_hits_14;
  wire                PmpPlugin_iGuard_hits_15;
  wire                when_PmpPlugin_l299;
  wire       [15:0]   _zz_IBusCachedPlugin_mmuBus_rsp_allowExecute;
  wire       [15:0]   _zz_IBusCachedPlugin_mmuBus_rsp_allowExecute_1;
  wire                _zz_IBusCachedPlugin_mmuBus_rsp_allowExecute_2;
  wire                _zz_IBusCachedPlugin_mmuBus_rsp_allowExecute_3;
  wire                _zz_IBusCachedPlugin_mmuBus_rsp_allowExecute_4;
  wire                _zz_IBusCachedPlugin_mmuBus_rsp_allowExecute_5;
  wire                _zz_IBusCachedPlugin_mmuBus_rsp_allowExecute_6;
  wire                _zz_IBusCachedPlugin_mmuBus_rsp_allowExecute_7;
  wire                _zz_IBusCachedPlugin_mmuBus_rsp_allowExecute_8;
  wire                _zz_IBusCachedPlugin_mmuBus_rsp_allowExecute_9;
  wire                _zz_IBusCachedPlugin_mmuBus_rsp_allowExecute_10;
  wire                _zz_IBusCachedPlugin_mmuBus_rsp_allowExecute_11;
  wire                _zz_IBusCachedPlugin_mmuBus_rsp_allowExecute_12;
  wire                _zz_IBusCachedPlugin_mmuBus_rsp_allowExecute_13;
  wire                _zz_IBusCachedPlugin_mmuBus_rsp_allowExecute_14;
  wire                _zz_IBusCachedPlugin_mmuBus_rsp_allowExecute_15;
  wire                _zz_IBusCachedPlugin_mmuBus_rsp_allowExecute_16;
  wire       [31:0]   _zz_decode_IS_RS2_SIGNED;
  wire                _zz_decode_IS_RS2_SIGNED_1;
  wire                _zz_decode_IS_RS2_SIGNED_2;
  wire                _zz_decode_IS_RS2_SIGNED_3;
  wire                _zz_decode_IS_RS2_SIGNED_4;
  wire                _zz_decode_IS_RS2_SIGNED_5;
  wire       [1:0]    _zz_decode_SRC1_CTRL_2;
  wire       [1:0]    _zz_decode_ALU_CTRL_2;
  wire       [1:0]    _zz_decode_SRC2_CTRL_2;
  wire       [1:0]    _zz_decode_ALU_BITWISE_CTRL_2;
  wire       [1:0]    _zz_decode_SHIFT_CTRL_2;
  wire       [1:0]    _zz_decode_BRANCH_CTRL_2;
  wire       [1:0]    _zz_decode_ENV_CTRL_2;
  wire                when_RegFilePlugin_l63;
  wire       [4:0]    decode_RegFilePlugin_regFileReadAddress1;
  wire       [4:0]    decode_RegFilePlugin_regFileReadAddress2;
  wire       [31:0]   decode_RegFilePlugin_rs1Data;
  wire       [31:0]   decode_RegFilePlugin_rs2Data;
  reg                 lastStageRegFileWrite_valid /* verilator public */ ;
  reg        [4:0]    lastStageRegFileWrite_payload_address /* verilator public */ ;
  reg        [31:0]   lastStageRegFileWrite_payload_data /* verilator public */ ;
  reg                 _zz_10;
  reg        [31:0]   execute_IntAluPlugin_bitwise;
  reg        [31:0]   _zz_execute_REGFILE_WRITE_DATA;
  reg        [31:0]   _zz_execute_SRC1;
  wire                _zz_execute_SRC2_1;
  reg        [19:0]   _zz_execute_SRC2_2;
  wire                _zz_execute_SRC2_3;
  reg        [19:0]   _zz_execute_SRC2_4;
  reg        [31:0]   _zz_execute_SRC2_5;
  reg        [31:0]   execute_SrcPlugin_addSub;
  wire                execute_SrcPlugin_less;
  wire       [4:0]    execute_FullBarrelShifterPlugin_amplitude;
  reg        [31:0]   _zz_execute_FullBarrelShifterPlugin_reversed;
  wire       [31:0]   execute_FullBarrelShifterPlugin_reversed;
  reg        [31:0]   _zz_decode_RS2_3;
  reg                 HazardSimplePlugin_src0Hazard;
  reg                 HazardSimplePlugin_src1Hazard;
  wire                HazardSimplePlugin_writeBackWrites_valid;
  wire       [4:0]    HazardSimplePlugin_writeBackWrites_payload_address;
  wire       [31:0]   HazardSimplePlugin_writeBackWrites_payload_data;
  reg                 HazardSimplePlugin_writeBackBuffer_valid;
  reg        [4:0]    HazardSimplePlugin_writeBackBuffer_payload_address;
  reg        [31:0]   HazardSimplePlugin_writeBackBuffer_payload_data;
  wire                HazardSimplePlugin_addr0Match;
  wire                HazardSimplePlugin_addr1Match;
  wire                when_HazardSimplePlugin_l47;
  wire                when_HazardSimplePlugin_l48;
  wire                when_HazardSimplePlugin_l51;
  wire                when_HazardSimplePlugin_l45;
  wire                when_HazardSimplePlugin_l57;
  wire                when_HazardSimplePlugin_l58;
  wire                when_HazardSimplePlugin_l48_1;
  wire                when_HazardSimplePlugin_l51_1;
  wire                when_HazardSimplePlugin_l45_1;
  wire                when_HazardSimplePlugin_l57_1;
  wire                when_HazardSimplePlugin_l58_1;
  wire                when_HazardSimplePlugin_l48_2;
  wire                when_HazardSimplePlugin_l51_2;
  wire                when_HazardSimplePlugin_l45_2;
  wire                when_HazardSimplePlugin_l57_2;
  wire                when_HazardSimplePlugin_l58_2;
  wire                when_HazardSimplePlugin_l105;
  wire                when_HazardSimplePlugin_l108;
  wire                when_HazardSimplePlugin_l113;
  wire                execute_BranchPlugin_eq;
  wire       [2:0]    switch_Misc_l210_1;
  reg                 _zz_execute_BRANCH_COND_RESULT;
  reg                 _zz_execute_BRANCH_COND_RESULT_1;
  wire                _zz_execute_BranchPlugin_missAlignedTarget;
  reg        [19:0]   _zz_execute_BranchPlugin_missAlignedTarget_1;
  wire                _zz_execute_BranchPlugin_missAlignedTarget_2;
  reg        [10:0]   _zz_execute_BranchPlugin_missAlignedTarget_3;
  wire                _zz_execute_BranchPlugin_missAlignedTarget_4;
  reg        [18:0]   _zz_execute_BranchPlugin_missAlignedTarget_5;
  reg                 _zz_execute_BranchPlugin_missAlignedTarget_6;
  wire                execute_BranchPlugin_missAlignedTarget;
  reg        [31:0]   execute_BranchPlugin_branch_src1;
  reg        [31:0]   execute_BranchPlugin_branch_src2;
  wire                _zz_execute_BranchPlugin_branch_src2;
  reg        [19:0]   _zz_execute_BranchPlugin_branch_src2_1;
  wire                _zz_execute_BranchPlugin_branch_src2_2;
  reg        [10:0]   _zz_execute_BranchPlugin_branch_src2_3;
  wire                _zz_execute_BranchPlugin_branch_src2_4;
  reg        [18:0]   _zz_execute_BranchPlugin_branch_src2_5;
  wire       [31:0]   execute_BranchPlugin_branchAdder;
  reg        [1:0]    _zz_CsrPlugin_privilege;
  reg        [1:0]    CsrPlugin_misa_base;
  reg        [25:0]   CsrPlugin_misa_extensions;
  reg        [1:0]    CsrPlugin_mtvec_mode;
  reg        [29:0]   CsrPlugin_mtvec_base;
  reg        [31:0]   CsrPlugin_mepc;
  reg                 CsrPlugin_mstatus_MIE;
  reg                 CsrPlugin_mstatus_MPIE;
  reg        [1:0]    CsrPlugin_mstatus_MPP;
  reg                 CsrPlugin_mip_MEIP;
  reg                 CsrPlugin_mip_MTIP;
  reg                 CsrPlugin_mip_MSIP;
  reg                 CsrPlugin_mie_MEIE;
  reg                 CsrPlugin_mie_MTIE;
  reg                 CsrPlugin_mie_MSIE;
  reg        [31:0]   CsrPlugin_mscratch;
  reg                 CsrPlugin_mcause_interrupt;
  reg        [3:0]    CsrPlugin_mcause_exceptionCode;
  reg        [31:0]   CsrPlugin_mtval;
  reg        [63:0]   CsrPlugin_mcycle;
  reg        [63:0]   CsrPlugin_minstret;
  wire                _zz_when_CsrPlugin_l965;
  wire                _zz_when_CsrPlugin_l965_1;
  wire                _zz_when_CsrPlugin_l965_2;
  reg                 CsrPlugin_exceptionPortCtrl_exceptionValids_decode;
  reg                 CsrPlugin_exceptionPortCtrl_exceptionValids_execute;
  reg                 CsrPlugin_exceptionPortCtrl_exceptionValids_memory;
  reg                 CsrPlugin_exceptionPortCtrl_exceptionValids_writeBack;
  reg                 CsrPlugin_exceptionPortCtrl_exceptionValidsRegs_decode;
  reg                 CsrPlugin_exceptionPortCtrl_exceptionValidsRegs_execute;
  reg                 CsrPlugin_exceptionPortCtrl_exceptionValidsRegs_memory;
  reg                 CsrPlugin_exceptionPortCtrl_exceptionValidsRegs_writeBack;
  reg        [3:0]    CsrPlugin_exceptionPortCtrl_exceptionContext_code;
  reg        [31:0]   CsrPlugin_exceptionPortCtrl_exceptionContext_badAddr;
  wire       [1:0]    CsrPlugin_exceptionPortCtrl_exceptionTargetPrivilegeUncapped;
  wire       [1:0]    CsrPlugin_exceptionPortCtrl_exceptionTargetPrivilege;
  wire       [1:0]    _zz_CsrPlugin_exceptionPortCtrl_exceptionContext_code;
  wire                _zz_CsrPlugin_exceptionPortCtrl_exceptionContext_code_1;
  wire                when_CsrPlugin_l922;
  wire                when_CsrPlugin_l922_1;
  wire                when_CsrPlugin_l922_2;
  wire                when_CsrPlugin_l922_3;
  wire                when_CsrPlugin_l935;
  reg                 CsrPlugin_interrupt_valid;
  reg        [3:0]    CsrPlugin_interrupt_code /* verilator public */ ;
  reg        [1:0]    CsrPlugin_interrupt_targetPrivilege;
  wire                when_CsrPlugin_l959;
  wire                when_CsrPlugin_l965;
  wire                when_CsrPlugin_l965_1;
  wire                when_CsrPlugin_l965_2;
  wire                CsrPlugin_exception;
  reg                 CsrPlugin_lastStageWasWfi;
  reg                 CsrPlugin_pipelineLiberator_pcValids_0;
  reg                 CsrPlugin_pipelineLiberator_pcValids_1;
  reg                 CsrPlugin_pipelineLiberator_pcValids_2;
  wire                CsrPlugin_pipelineLiberator_active;
  wire                when_CsrPlugin_l993;
  wire                when_CsrPlugin_l993_1;
  wire                when_CsrPlugin_l993_2;
  wire                when_CsrPlugin_l998;
  reg                 CsrPlugin_pipelineLiberator_done;
  wire                when_CsrPlugin_l1004;
  wire                CsrPlugin_interruptJump /* verilator public */ ;
  reg                 CsrPlugin_hadException /* verilator public */ ;
  reg        [1:0]    CsrPlugin_targetPrivilege;
  reg        [3:0]    CsrPlugin_trapCause;
  reg        [1:0]    CsrPlugin_xtvec_mode;
  reg        [29:0]   CsrPlugin_xtvec_base;
  wire                when_CsrPlugin_l1032;
  wire                when_CsrPlugin_l1077;
  wire       [1:0]    switch_CsrPlugin_l1081;
  reg                 execute_CsrPlugin_wfiWake;
  wire                when_CsrPlugin_l1121;
  wire                when_CsrPlugin_l1123;
  wire                when_CsrPlugin_l1129;
  wire                execute_CsrPlugin_blockedBySideEffects;
  reg                 execute_CsrPlugin_illegalAccess;
  reg                 execute_CsrPlugin_illegalInstruction;
  wire                when_CsrPlugin_l1142;
  wire                when_CsrPlugin_l1149;
  wire                when_CsrPlugin_l1150;
  wire                when_CsrPlugin_l1157;
  reg                 execute_CsrPlugin_writeInstruction;
  reg                 execute_CsrPlugin_readInstruction;
  wire                execute_CsrPlugin_writeEnable;
  wire                execute_CsrPlugin_readEnable;
  wire       [31:0]   execute_CsrPlugin_readToWriteData;
  wire                switch_Misc_l210_2;
  reg        [31:0]   _zz_CsrPlugin_csrMapping_writeDataSignal;
  wire                when_CsrPlugin_l1189;
  wire                when_CsrPlugin_l1193;
  wire       [11:0]   execute_CsrPlugin_csrAddress;
  reg                 execute_MulPlugin_aSigned;
  reg                 execute_MulPlugin_bSigned;
  wire       [31:0]   execute_MulPlugin_a;
  wire       [31:0]   execute_MulPlugin_b;
  wire       [1:0]    switch_MulPlugin_l87;
  wire       [15:0]   execute_MulPlugin_aULow;
  wire       [15:0]   execute_MulPlugin_bULow;
  wire       [16:0]   execute_MulPlugin_aSLow;
  wire       [16:0]   execute_MulPlugin_bSLow;
  wire       [16:0]   execute_MulPlugin_aHigh;
  wire       [16:0]   execute_MulPlugin_bHigh;
  wire       [65:0]   writeBack_MulPlugin_result;
  wire                when_MulPlugin_l147;
  wire       [1:0]    switch_MulPlugin_l148;
  reg        [32:0]   memory_DivPlugin_rs1;
  reg        [31:0]   memory_DivPlugin_rs2;
  reg        [64:0]   memory_DivPlugin_accumulator;
  wire                memory_DivPlugin_frontendOk;
  reg                 memory_DivPlugin_div_needRevert;
  reg                 memory_DivPlugin_div_counter_willIncrement;
  reg                 memory_DivPlugin_div_counter_willClear;
  reg        [5:0]    memory_DivPlugin_div_counter_valueNext;
  reg        [5:0]    memory_DivPlugin_div_counter_value;
  wire                memory_DivPlugin_div_counter_willOverflowIfInc;
  wire                memory_DivPlugin_div_counter_willOverflow;
  reg                 memory_DivPlugin_div_done;
  wire                when_MulDivIterativePlugin_l126;
  wire                when_MulDivIterativePlugin_l126_1;
  reg        [31:0]   memory_DivPlugin_div_result;
  wire                when_MulDivIterativePlugin_l128;
  wire                when_MulDivIterativePlugin_l129;
  wire                when_MulDivIterativePlugin_l132;
  wire       [31:0]   _zz_memory_DivPlugin_div_stage_0_remainderShifted;
  wire       [32:0]   memory_DivPlugin_div_stage_0_remainderShifted;
  wire       [32:0]   memory_DivPlugin_div_stage_0_remainderMinusDenominator;
  wire       [31:0]   memory_DivPlugin_div_stage_0_outRemainder;
  wire       [31:0]   memory_DivPlugin_div_stage_0_outNumerator;
  wire                when_MulDivIterativePlugin_l151;
  wire       [31:0]   _zz_memory_DivPlugin_div_result;
  wire                when_MulDivIterativePlugin_l162;
  wire                _zz_memory_DivPlugin_rs2;
  wire                _zz_memory_DivPlugin_rs1;
  reg        [32:0]   _zz_memory_DivPlugin_rs1_1;
  reg        [31:0]   externalInterruptArray_regNext;
  reg        [31:0]   _zz_CsrPlugin_csrMapping_readDataInit;
  wire       [31:0]   _zz_CsrPlugin_csrMapping_readDataInit_1;
  wire                when_Pipeline_l124;
  reg        [31:0]   decode_to_execute_PC;
  wire                when_Pipeline_l124_1;
  reg        [31:0]   execute_to_memory_PC;
  wire                when_Pipeline_l124_2;
  reg        [31:0]   memory_to_writeBack_PC;
  wire                when_Pipeline_l124_3;
  reg        [31:0]   decode_to_execute_INSTRUCTION;
  wire                when_Pipeline_l124_4;
  reg        [31:0]   execute_to_memory_INSTRUCTION;
  wire                when_Pipeline_l124_5;
  reg        [31:0]   memory_to_writeBack_INSTRUCTION;
  wire                when_Pipeline_l124_6;
  reg        [31:0]   decode_to_execute_FORMAL_PC_NEXT;
  wire                when_Pipeline_l124_7;
  reg        [31:0]   execute_to_memory_FORMAL_PC_NEXT;
  wire                when_Pipeline_l124_8;
  reg        [31:0]   memory_to_writeBack_FORMAL_PC_NEXT;
  wire                when_Pipeline_l124_9;
  reg                 decode_to_execute_MEMORY_FORCE_CONSTISTENCY;
  wire                when_Pipeline_l124_10;
  reg        [1:0]    decode_to_execute_SRC1_CTRL;
  wire                when_Pipeline_l124_11;
  reg                 decode_to_execute_SRC_USE_SUB_LESS;
  wire                when_Pipeline_l124_12;
  reg                 decode_to_execute_MEMORY_ENABLE;
  wire                when_Pipeline_l124_13;
  reg                 execute_to_memory_MEMORY_ENABLE;
  wire                when_Pipeline_l124_14;
  reg                 memory_to_writeBack_MEMORY_ENABLE;
  wire                when_Pipeline_l124_15;
  reg        [1:0]    decode_to_execute_ALU_CTRL;
  wire                when_Pipeline_l124_16;
  reg        [1:0]    decode_to_execute_SRC2_CTRL;
  wire                when_Pipeline_l124_17;
  reg                 decode_to_execute_REGFILE_WRITE_VALID;
  wire                when_Pipeline_l124_18;
  reg                 execute_to_memory_REGFILE_WRITE_VALID;
  wire                when_Pipeline_l124_19;
  reg                 memory_to_writeBack_REGFILE_WRITE_VALID;
  wire                when_Pipeline_l124_20;
  reg                 decode_to_execute_BYPASSABLE_EXECUTE_STAGE;
  wire                when_Pipeline_l124_21;
  reg                 decode_to_execute_BYPASSABLE_MEMORY_STAGE;
  wire                when_Pipeline_l124_22;
  reg                 execute_to_memory_BYPASSABLE_MEMORY_STAGE;
  wire                when_Pipeline_l124_23;
  reg                 decode_to_execute_MEMORY_WR;
  wire                when_Pipeline_l124_24;
  reg                 execute_to_memory_MEMORY_WR;
  wire                when_Pipeline_l124_25;
  reg                 memory_to_writeBack_MEMORY_WR;
  wire                when_Pipeline_l124_26;
  reg                 decode_to_execute_MEMORY_MANAGMENT;
  wire                when_Pipeline_l124_27;
  reg                 decode_to_execute_SRC_LESS_UNSIGNED;
  wire                when_Pipeline_l124_28;
  reg        [1:0]    decode_to_execute_ALU_BITWISE_CTRL;
  wire                when_Pipeline_l124_29;
  reg        [1:0]    decode_to_execute_SHIFT_CTRL;
  wire                when_Pipeline_l124_30;
  reg        [1:0]    execute_to_memory_SHIFT_CTRL;
  wire                when_Pipeline_l124_31;
  reg        [1:0]    decode_to_execute_BRANCH_CTRL;
  wire                when_Pipeline_l124_32;
  reg                 decode_to_execute_IS_CSR;
  wire                when_Pipeline_l124_33;
  reg        [1:0]    decode_to_execute_ENV_CTRL;
  wire                when_Pipeline_l124_34;
  reg        [1:0]    execute_to_memory_ENV_CTRL;
  wire                when_Pipeline_l124_35;
  reg        [1:0]    memory_to_writeBack_ENV_CTRL;
  wire                when_Pipeline_l124_36;
  reg                 decode_to_execute_IS_MUL;
  wire                when_Pipeline_l124_37;
  reg                 execute_to_memory_IS_MUL;
  wire                when_Pipeline_l124_38;
  reg                 memory_to_writeBack_IS_MUL;
  wire                when_Pipeline_l124_39;
  reg                 decode_to_execute_IS_DIV;
  wire                when_Pipeline_l124_40;
  reg                 execute_to_memory_IS_DIV;
  wire                when_Pipeline_l124_41;
  reg                 decode_to_execute_IS_RS1_SIGNED;
  wire                when_Pipeline_l124_42;
  reg                 decode_to_execute_IS_RS2_SIGNED;
  wire                when_Pipeline_l124_43;
  reg        [31:0]   decode_to_execute_RS1;
  wire                when_Pipeline_l124_44;
  reg        [31:0]   decode_to_execute_RS2;
  wire                when_Pipeline_l124_45;
  reg                 decode_to_execute_SRC2_FORCE_ZERO;
  wire                when_Pipeline_l124_46;
  reg                 decode_to_execute_PREDICTION_HAD_BRANCHED2;
  wire                when_Pipeline_l124_47;
  reg                 decode_to_execute_CSR_WRITE_OPCODE;
  wire                when_Pipeline_l124_48;
  reg                 decode_to_execute_CSR_READ_OPCODE;
  wire                when_Pipeline_l124_49;
  reg        [31:0]   execute_to_memory_MEMORY_STORE_DATA_RF;
  wire                when_Pipeline_l124_50;
  reg        [31:0]   memory_to_writeBack_MEMORY_STORE_DATA_RF;
  wire                when_Pipeline_l124_51;
  reg        [31:0]   execute_to_memory_REGFILE_WRITE_DATA;
  wire                when_Pipeline_l124_52;
  reg        [31:0]   memory_to_writeBack_REGFILE_WRITE_DATA;
  wire                when_Pipeline_l124_53;
  reg        [31:0]   execute_to_memory_SHIFT_RIGHT;
  wire                when_Pipeline_l124_54;
  reg                 execute_to_memory_BRANCH_DO;
  wire                when_Pipeline_l124_55;
  reg        [31:0]   execute_to_memory_BRANCH_CALC;
  wire                when_Pipeline_l124_56;
  reg        [31:0]   execute_to_memory_MUL_LL;
  wire                when_Pipeline_l124_57;
  reg        [33:0]   execute_to_memory_MUL_LH;
  wire                when_Pipeline_l124_58;
  reg        [33:0]   execute_to_memory_MUL_HL;
  wire                when_Pipeline_l124_59;
  reg        [33:0]   execute_to_memory_MUL_HH;
  wire                when_Pipeline_l124_60;
  reg        [33:0]   memory_to_writeBack_MUL_HH;
  wire                when_Pipeline_l124_61;
  reg        [51:0]   memory_to_writeBack_MUL_LOW;
  wire                when_Pipeline_l151;
  wire                when_Pipeline_l154;
  wire                when_Pipeline_l151_1;
  wire                when_Pipeline_l154_1;
  wire                when_Pipeline_l151_2;
  wire                when_Pipeline_l154_2;
  reg        [2:0]    execute_PmpPlugin_fsm_stateReg;
  reg        [2:0]    execute_PmpPlugin_fsm_stateNext;
  wire       [7:0]    _zz_PmpPlugin_pmpcfg_0;
  wire       [7:0]    _zz_PmpPlugin_pmpcfg_0_1;
  wire       [7:0]    _zz_PmpPlugin_pmpcfg_0_2;
  wire       [7:0]    _zz_PmpPlugin_pmpcfg_0_3;
  wire                when_PmpPlugin_l209;
  wire       [15:0]   _zz_11;
  wire                when_PmpPlugin_l209_1;
  wire       [15:0]   _zz_12;
  wire                when_PmpPlugin_l209_2;
  wire       [15:0]   _zz_13;
  wire                when_PmpPlugin_l209_3;
  wire       [15:0]   _zz_14;
  wire                when_PmpPlugin_l216;
  wire                when_PmpPlugin_l229;
  wire                when_StateMachine_l233;
  wire                when_StateMachine_l249;
  wire                when_StateMachine_l249_1;
  wire                when_StateMachine_l249_2;
  wire                when_CsrPlugin_l1277;
  reg                 execute_CsrPlugin_csr_3264;
  wire                when_CsrPlugin_l1277_1;
  reg                 execute_CsrPlugin_csr_3857;
  wire                when_CsrPlugin_l1277_2;
  reg                 execute_CsrPlugin_csr_3858;
  wire                when_CsrPlugin_l1277_3;
  reg                 execute_CsrPlugin_csr_3859;
  wire                when_CsrPlugin_l1277_4;
  reg                 execute_CsrPlugin_csr_3860;
  wire                when_CsrPlugin_l1277_5;
  reg                 execute_CsrPlugin_csr_769;
  wire                when_CsrPlugin_l1277_6;
  reg                 execute_CsrPlugin_csr_768;
  wire                when_CsrPlugin_l1277_7;
  reg                 execute_CsrPlugin_csr_836;
  wire                when_CsrPlugin_l1277_8;
  reg                 execute_CsrPlugin_csr_772;
  wire                when_CsrPlugin_l1277_9;
  reg                 execute_CsrPlugin_csr_773;
  wire                when_CsrPlugin_l1277_10;
  reg                 execute_CsrPlugin_csr_833;
  wire                when_CsrPlugin_l1277_11;
  reg                 execute_CsrPlugin_csr_832;
  wire                when_CsrPlugin_l1277_12;
  reg                 execute_CsrPlugin_csr_834;
  wire                when_CsrPlugin_l1277_13;
  reg                 execute_CsrPlugin_csr_835;
  wire                when_CsrPlugin_l1277_14;
  reg                 execute_CsrPlugin_csr_2816;
  wire                when_CsrPlugin_l1277_15;
  reg                 execute_CsrPlugin_csr_2944;
  wire                when_CsrPlugin_l1277_16;
  reg                 execute_CsrPlugin_csr_2818;
  wire                when_CsrPlugin_l1277_17;
  reg                 execute_CsrPlugin_csr_2946;
  wire                when_CsrPlugin_l1277_18;
  reg                 execute_CsrPlugin_csr_3072;
  wire                when_CsrPlugin_l1277_19;
  reg                 execute_CsrPlugin_csr_3200;
  wire                when_CsrPlugin_l1277_20;
  reg                 execute_CsrPlugin_csr_3074;
  wire                when_CsrPlugin_l1277_21;
  reg                 execute_CsrPlugin_csr_3202;
  wire                when_CsrPlugin_l1277_22;
  reg                 execute_CsrPlugin_csr_3008;
  wire                when_CsrPlugin_l1277_23;
  reg                 execute_CsrPlugin_csr_4032;
  reg        [31:0]   _zz_CsrPlugin_csrMapping_readDataInit_2;
  reg        [31:0]   _zz_CsrPlugin_csrMapping_readDataInit_3;
  reg        [31:0]   _zz_CsrPlugin_csrMapping_readDataInit_4;
  reg        [31:0]   _zz_CsrPlugin_csrMapping_readDataInit_5;
  reg        [31:0]   _zz_CsrPlugin_csrMapping_readDataInit_6;
  wire       [1:0]    switch_CsrPlugin_l723;
  reg        [31:0]   _zz_CsrPlugin_csrMapping_readDataInit_7;
  reg        [31:0]   _zz_CsrPlugin_csrMapping_readDataInit_8;
  reg        [31:0]   _zz_CsrPlugin_csrMapping_readDataInit_9;
  reg        [31:0]   _zz_CsrPlugin_csrMapping_readDataInit_10;
  reg        [31:0]   _zz_CsrPlugin_csrMapping_readDataInit_11;
  reg        [31:0]   _zz_CsrPlugin_csrMapping_readDataInit_12;
  reg        [31:0]   _zz_CsrPlugin_csrMapping_readDataInit_13;
  reg        [31:0]   _zz_CsrPlugin_csrMapping_readDataInit_14;
  reg        [31:0]   _zz_CsrPlugin_csrMapping_readDataInit_15;
  reg        [31:0]   _zz_CsrPlugin_csrMapping_readDataInit_16;
  reg        [31:0]   _zz_CsrPlugin_csrMapping_readDataInit_17;
  reg        [31:0]   _zz_CsrPlugin_csrMapping_readDataInit_18;
  reg        [31:0]   _zz_CsrPlugin_csrMapping_readDataInit_19;
  reg        [31:0]   _zz_CsrPlugin_csrMapping_readDataInit_20;
  reg        [31:0]   _zz_CsrPlugin_csrMapping_readDataInit_21;
  reg        [31:0]   _zz_CsrPlugin_csrMapping_readDataInit_22;
  reg        [31:0]   _zz_CsrPlugin_csrMapping_readDataInit_23;
  reg        [31:0]   _zz_CsrPlugin_csrMapping_readDataInit_24;
  wire                when_PmpPlugin_l155;
  wire                when_PmpPlugin_l172;
  wire                when_PmpPlugin_l175;
  wire                when_CsrPlugin_l1310;
  wire                when_CsrPlugin_l1315;
  reg        [2:0]    _zz_iBusWishbone_ADR;
  wire                when_InstructionCache_l239;
  reg                 _zz_iBus_rsp_valid;
  reg        [31:0]   iBusWishbone_DAT_MISO_regNext;
  reg        [2:0]    _zz_dBus_cmd_ready;
  wire                _zz_dBus_cmd_ready_1;
  wire                _zz_dBus_cmd_ready_2;
  wire                _zz_dBus_cmd_ready_3;
  wire                _zz_dBus_cmd_ready_4;
  wire                _zz_dBus_cmd_ready_5;
  reg                 _zz_dBus_rsp_valid;
  reg        [31:0]   dBusWishbone_DAT_MISO_regNext;
  `ifndef SYNTHESIS
  reg [39:0] _zz_memory_to_writeBack_ENV_CTRL_string;
  reg [39:0] _zz_memory_to_writeBack_ENV_CTRL_1_string;
  reg [39:0] _zz_execute_to_memory_ENV_CTRL_string;
  reg [39:0] _zz_execute_to_memory_ENV_CTRL_1_string;
  reg [39:0] decode_ENV_CTRL_string;
  reg [39:0] _zz_decode_ENV_CTRL_string;
  reg [39:0] _zz_decode_to_execute_ENV_CTRL_string;
  reg [39:0] _zz_decode_to_execute_ENV_CTRL_1_string;
  reg [31:0] _zz_decode_to_execute_BRANCH_CTRL_string;
  reg [31:0] _zz_decode_to_execute_BRANCH_CTRL_1_string;
  reg [71:0] _zz_execute_to_memory_SHIFT_CTRL_string;
  reg [71:0] _zz_execute_to_memory_SHIFT_CTRL_1_string;
  reg [71:0] decode_SHIFT_CTRL_string;
  reg [71:0] _zz_decode_SHIFT_CTRL_string;
  reg [71:0] _zz_decode_to_execute_SHIFT_CTRL_string;
  reg [71:0] _zz_decode_to_execute_SHIFT_CTRL_1_string;
  reg [39:0] decode_ALU_BITWISE_CTRL_string;
  reg [39:0] _zz_decode_ALU_BITWISE_CTRL_string;
  reg [39:0] _zz_decode_to_execute_ALU_BITWISE_CTRL_string;
  reg [39:0] _zz_decode_to_execute_ALU_BITWISE_CTRL_1_string;
  reg [23:0] decode_SRC2_CTRL_string;
  reg [23:0] _zz_decode_SRC2_CTRL_string;
  reg [23:0] _zz_decode_to_execute_SRC2_CTRL_string;
  reg [23:0] _zz_decode_to_execute_SRC2_CTRL_1_string;
  reg [63:0] decode_ALU_CTRL_string;
  reg [63:0] _zz_decode_ALU_CTRL_string;
  reg [63:0] _zz_decode_to_execute_ALU_CTRL_string;
  reg [63:0] _zz_decode_to_execute_ALU_CTRL_1_string;
  reg [95:0] decode_SRC1_CTRL_string;
  reg [95:0] _zz_decode_SRC1_CTRL_string;
  reg [95:0] _zz_decode_to_execute_SRC1_CTRL_string;
  reg [95:0] _zz_decode_to_execute_SRC1_CTRL_1_string;
  reg [39:0] memory_ENV_CTRL_string;
  reg [39:0] _zz_memory_ENV_CTRL_string;
  reg [39:0] execute_ENV_CTRL_string;
  reg [39:0] _zz_execute_ENV_CTRL_string;
  reg [39:0] writeBack_ENV_CTRL_string;
  reg [39:0] _zz_writeBack_ENV_CTRL_string;
  reg [31:0] execute_BRANCH_CTRL_string;
  reg [31:0] _zz_execute_BRANCH_CTRL_string;
  reg [71:0] memory_SHIFT_CTRL_string;
  reg [71:0] _zz_memory_SHIFT_CTRL_string;
  reg [71:0] execute_SHIFT_CTRL_string;
  reg [71:0] _zz_execute_SHIFT_CTRL_string;
  reg [23:0] execute_SRC2_CTRL_string;
  reg [23:0] _zz_execute_SRC2_CTRL_string;
  reg [95:0] execute_SRC1_CTRL_string;
  reg [95:0] _zz_execute_SRC1_CTRL_string;
  reg [63:0] execute_ALU_CTRL_string;
  reg [63:0] _zz_execute_ALU_CTRL_string;
  reg [39:0] execute_ALU_BITWISE_CTRL_string;
  reg [39:0] _zz_execute_ALU_BITWISE_CTRL_string;
  reg [39:0] _zz_decode_ENV_CTRL_1_string;
  reg [31:0] _zz_decode_BRANCH_CTRL_string;
  reg [71:0] _zz_decode_SHIFT_CTRL_1_string;
  reg [39:0] _zz_decode_ALU_BITWISE_CTRL_1_string;
  reg [23:0] _zz_decode_SRC2_CTRL_1_string;
  reg [63:0] _zz_decode_ALU_CTRL_1_string;
  reg [95:0] _zz_decode_SRC1_CTRL_1_string;
  reg [31:0] decode_BRANCH_CTRL_string;
  reg [31:0] _zz_decode_BRANCH_CTRL_1_string;
  reg [95:0] _zz_decode_SRC1_CTRL_2_string;
  reg [63:0] _zz_decode_ALU_CTRL_2_string;
  reg [23:0] _zz_decode_SRC2_CTRL_2_string;
  reg [39:0] _zz_decode_ALU_BITWISE_CTRL_2_string;
  reg [71:0] _zz_decode_SHIFT_CTRL_2_string;
  reg [31:0] _zz_decode_BRANCH_CTRL_2_string;
  reg [39:0] _zz_decode_ENV_CTRL_2_string;
  reg [95:0] decode_to_execute_SRC1_CTRL_string;
  reg [63:0] decode_to_execute_ALU_CTRL_string;
  reg [23:0] decode_to_execute_SRC2_CTRL_string;
  reg [39:0] decode_to_execute_ALU_BITWISE_CTRL_string;
  reg [71:0] decode_to_execute_SHIFT_CTRL_string;
  reg [71:0] execute_to_memory_SHIFT_CTRL_string;
  reg [31:0] decode_to_execute_BRANCH_CTRL_string;
  reg [39:0] decode_to_execute_ENV_CTRL_string;
  reg [39:0] execute_to_memory_ENV_CTRL_string;
  reg [39:0] memory_to_writeBack_ENV_CTRL_string;
  reg [79:0] execute_PmpPlugin_fsm_stateReg_string;
  reg [79:0] execute_PmpPlugin_fsm_stateNext_string;
  `endif

  (* ram_style = "distributed" *) reg [31:0] PmpPlugin_pmpaddr [0:15];
  (* no_rw_check , ram_style = "block" *) reg [31:0] RegFilePlugin_regFile [0:31] /* verilator public */ ;

  assign _zz_when = ({decodeExceptionPort_valid,IBusCachedPlugin_decodeExceptionPort_valid} != 2'b00);
  assign _zz_memory_MUL_LOW = ($signed(_zz_memory_MUL_LOW_1) + $signed(_zz_memory_MUL_LOW_5));
  assign _zz_memory_MUL_LOW_1 = ($signed(_zz_memory_MUL_LOW_2) + $signed(_zz_memory_MUL_LOW_3));
  assign _zz_memory_MUL_LOW_2 = 52'h0;
  assign _zz_memory_MUL_LOW_4 = {1'b0,memory_MUL_LL};
  assign _zz_memory_MUL_LOW_3 = {{19{_zz_memory_MUL_LOW_4[32]}}, _zz_memory_MUL_LOW_4};
  assign _zz_memory_MUL_LOW_6 = ({16'd0,memory_MUL_LH} <<< 16);
  assign _zz_memory_MUL_LOW_5 = {{2{_zz_memory_MUL_LOW_6[49]}}, _zz_memory_MUL_LOW_6};
  assign _zz_memory_MUL_LOW_8 = ({16'd0,memory_MUL_HL} <<< 16);
  assign _zz_memory_MUL_LOW_7 = {{2{_zz_memory_MUL_LOW_8[49]}}, _zz_memory_MUL_LOW_8};
  assign _zz_execute_SHIFT_RIGHT_1 = ($signed(_zz_execute_SHIFT_RIGHT_2) >>> execute_FullBarrelShifterPlugin_amplitude);
  assign _zz_execute_SHIFT_RIGHT = _zz_execute_SHIFT_RIGHT_1[31 : 0];
  assign _zz_execute_SHIFT_RIGHT_2 = {((execute_SHIFT_CTRL == ShiftCtrlEnum_SRA_1) && execute_FullBarrelShifterPlugin_reversed[31]),execute_FullBarrelShifterPlugin_reversed};
  assign _zz__zz_IBusCachedPlugin_jump_pcLoad_payload_1 = (_zz_IBusCachedPlugin_jump_pcLoad_payload - 4'b0001);
  assign _zz_IBusCachedPlugin_fetchPc_pc_1 = {IBusCachedPlugin_fetchPc_inc,2'b00};
  assign _zz_IBusCachedPlugin_fetchPc_pc = {29'd0, _zz_IBusCachedPlugin_fetchPc_pc_1};
  assign _zz__zz_IBusCachedPlugin_decodePrediction_cmd_hadBranch = {{{decode_INSTRUCTION[31],decode_INSTRUCTION[7]},decode_INSTRUCTION[30 : 25]},decode_INSTRUCTION[11 : 8]};
  assign _zz_IBusCachedPlugin_decodePrediction_cmd_hadBranch_2 = {{_zz_IBusCachedPlugin_decodePrediction_cmd_hadBranch_1,{{{decode_INSTRUCTION[31],decode_INSTRUCTION[7]},decode_INSTRUCTION[30 : 25]},decode_INSTRUCTION[11 : 8]}},1'b0};
  assign _zz__zz_3 = {{{decode_INSTRUCTION[31],decode_INSTRUCTION[19 : 12]},decode_INSTRUCTION[20]},decode_INSTRUCTION[30 : 21]};
  assign _zz__zz_5 = {{{decode_INSTRUCTION[31],decode_INSTRUCTION[7]},decode_INSTRUCTION[30 : 25]},decode_INSTRUCTION[11 : 8]};
  assign _zz__zz_7 = {{_zz_4,{{{decode_INSTRUCTION[31],decode_INSTRUCTION[19 : 12]},decode_INSTRUCTION[20]},decode_INSTRUCTION[30 : 21]}},1'b0};
  assign _zz__zz_7_1 = {{_zz_6,{{{decode_INSTRUCTION[31],decode_INSTRUCTION[7]},decode_INSTRUCTION[30 : 25]},decode_INSTRUCTION[11 : 8]}},1'b0};
  assign _zz__zz_IBusCachedPlugin_predictionJumpInterface_payload = {{{decode_INSTRUCTION[31],decode_INSTRUCTION[19 : 12]},decode_INSTRUCTION[20]},decode_INSTRUCTION[30 : 21]};
  assign _zz__zz_IBusCachedPlugin_predictionJumpInterface_payload_2 = {{{decode_INSTRUCTION[31],decode_INSTRUCTION[7]},decode_INSTRUCTION[30 : 25]},decode_INSTRUCTION[11 : 8]};
  assign _zz_io_cpu_flush_payload_lineId = _zz_io_cpu_flush_payload_lineId_1;
  assign _zz_io_cpu_flush_payload_lineId_1 = (execute_RS1 >>> 5);
  assign _zz_DBusCachedPlugin_exceptionBus_payload_code = (writeBack_MEMORY_WR ? 3'b111 : 3'b101);
  assign _zz_DBusCachedPlugin_exceptionBus_payload_code_1 = (writeBack_MEMORY_WR ? 3'b110 : 3'b100);
  assign _zz__zz_DBusCachedPlugin_mmuBus_rsp_allowRead_1_1 = (_zz_DBusCachedPlugin_mmuBus_rsp_allowRead - 16'h0001);
  assign _zz__zz_DBusCachedPlugin_mmuBus_rsp_allowWrite_1_1 = (_zz_DBusCachedPlugin_mmuBus_rsp_allowWrite - 16'h0001);
  assign _zz__zz_IBusCachedPlugin_mmuBus_rsp_allowExecute_1_1 = (_zz_IBusCachedPlugin_mmuBus_rsp_allowExecute - 16'h0001);
  assign _zz__zz_execute_REGFILE_WRITE_DATA = execute_SRC_LESS;
  assign _zz__zz_execute_SRC1 = 3'b100;
  assign _zz__zz_execute_SRC1_1 = execute_INSTRUCTION[19 : 15];
  assign _zz__zz_execute_SRC2_3 = {execute_INSTRUCTION[31 : 25],execute_INSTRUCTION[11 : 7]};
  assign _zz_execute_SrcPlugin_addSub = ($signed(_zz_execute_SrcPlugin_addSub_1) + $signed(_zz_execute_SrcPlugin_addSub_4));
  assign _zz_execute_SrcPlugin_addSub_1 = ($signed(_zz_execute_SrcPlugin_addSub_2) + $signed(_zz_execute_SrcPlugin_addSub_3));
  assign _zz_execute_SrcPlugin_addSub_2 = execute_SRC1;
  assign _zz_execute_SrcPlugin_addSub_3 = (execute_SRC_USE_SUB_LESS ? (~ execute_SRC2) : execute_SRC2);
  assign _zz_execute_SrcPlugin_addSub_4 = (execute_SRC_USE_SUB_LESS ? _zz_execute_SrcPlugin_addSub_5 : _zz_execute_SrcPlugin_addSub_6);
  assign _zz_execute_SrcPlugin_addSub_5 = 32'h00000001;
  assign _zz_execute_SrcPlugin_addSub_6 = 32'h0;
  assign _zz__zz_execute_BranchPlugin_missAlignedTarget_2 = {{{execute_INSTRUCTION[31],execute_INSTRUCTION[19 : 12]},execute_INSTRUCTION[20]},execute_INSTRUCTION[30 : 21]};
  assign _zz__zz_execute_BranchPlugin_missAlignedTarget_4 = {{{execute_INSTRUCTION[31],execute_INSTRUCTION[7]},execute_INSTRUCTION[30 : 25]},execute_INSTRUCTION[11 : 8]};
  assign _zz__zz_execute_BranchPlugin_missAlignedTarget_6 = {_zz_execute_BranchPlugin_missAlignedTarget_1,execute_INSTRUCTION[31 : 20]};
  assign _zz__zz_execute_BranchPlugin_missAlignedTarget_6_1 = {{_zz_execute_BranchPlugin_missAlignedTarget_3,{{{execute_INSTRUCTION[31],execute_INSTRUCTION[19 : 12]},execute_INSTRUCTION[20]},execute_INSTRUCTION[30 : 21]}},1'b0};
  assign _zz__zz_execute_BranchPlugin_missAlignedTarget_6_2 = {{_zz_execute_BranchPlugin_missAlignedTarget_5,{{{execute_INSTRUCTION[31],execute_INSTRUCTION[7]},execute_INSTRUCTION[30 : 25]},execute_INSTRUCTION[11 : 8]}},1'b0};
  assign _zz__zz_execute_BranchPlugin_branch_src2_2 = {{{execute_INSTRUCTION[31],execute_INSTRUCTION[19 : 12]},execute_INSTRUCTION[20]},execute_INSTRUCTION[30 : 21]};
  assign _zz__zz_execute_BranchPlugin_branch_src2_4 = {{{execute_INSTRUCTION[31],execute_INSTRUCTION[7]},execute_INSTRUCTION[30 : 25]},execute_INSTRUCTION[11 : 8]};
  assign _zz_execute_BranchPlugin_branch_src2_9 = 3'b100;
  assign _zz__zz_CsrPlugin_exceptionPortCtrl_exceptionContext_code_1 = (_zz_CsrPlugin_exceptionPortCtrl_exceptionContext_code & (~ _zz__zz_CsrPlugin_exceptionPortCtrl_exceptionContext_code_1_1));
  assign _zz__zz_CsrPlugin_exceptionPortCtrl_exceptionContext_code_1_1 = (_zz_CsrPlugin_exceptionPortCtrl_exceptionContext_code - 2'b01);
  assign _zz_writeBack_MulPlugin_result = {{14{writeBack_MUL_LOW[51]}}, writeBack_MUL_LOW};
  assign _zz_writeBack_MulPlugin_result_1 = ({32'd0,writeBack_MUL_HH} <<< 32);
  assign _zz__zz_decode_RS2_2 = writeBack_MUL_LOW[31 : 0];
  assign _zz__zz_decode_RS2_2_1 = writeBack_MulPlugin_result[63 : 32];
  assign _zz_memory_DivPlugin_div_counter_valueNext_1 = memory_DivPlugin_div_counter_willIncrement;
  assign _zz_memory_DivPlugin_div_counter_valueNext = {5'd0, _zz_memory_DivPlugin_div_counter_valueNext_1};
  assign _zz_memory_DivPlugin_div_stage_0_remainderMinusDenominator = {1'd0, memory_DivPlugin_rs2};
  assign _zz_memory_DivPlugin_div_stage_0_outRemainder = memory_DivPlugin_div_stage_0_remainderMinusDenominator[31:0];
  assign _zz_memory_DivPlugin_div_stage_0_outRemainder_1 = memory_DivPlugin_div_stage_0_remainderShifted[31:0];
  assign _zz_memory_DivPlugin_div_stage_0_outNumerator = {_zz_memory_DivPlugin_div_stage_0_remainderShifted,(! memory_DivPlugin_div_stage_0_remainderMinusDenominator[32])};
  assign _zz_memory_DivPlugin_div_result_1 = _zz_memory_DivPlugin_div_result_2;
  assign _zz_memory_DivPlugin_div_result_2 = _zz_memory_DivPlugin_div_result_3;
  assign _zz_memory_DivPlugin_div_result_3 = ({memory_DivPlugin_div_needRevert,(memory_DivPlugin_div_needRevert ? (~ _zz_memory_DivPlugin_div_result) : _zz_memory_DivPlugin_div_result)} + _zz_memory_DivPlugin_div_result_4);
  assign _zz_memory_DivPlugin_div_result_5 = memory_DivPlugin_div_needRevert;
  assign _zz_memory_DivPlugin_div_result_4 = {32'd0, _zz_memory_DivPlugin_div_result_5};
  assign _zz_memory_DivPlugin_rs1_3 = _zz_memory_DivPlugin_rs1;
  assign _zz_memory_DivPlugin_rs1_2 = {32'd0, _zz_memory_DivPlugin_rs1_3};
  assign _zz_memory_DivPlugin_rs2_2 = _zz_memory_DivPlugin_rs2;
  assign _zz_memory_DivPlugin_rs2_1 = {31'd0, _zz_memory_DivPlugin_rs2_2};
  assign _zz_iBusWishbone_ADR_1 = (iBus_cmd_payload_address >>> 5);
  assign _zz_PmpPlugin_pmpaddr_port = execute_PmpPlugin_writeData_;
  assign _zz_decode_RegFilePlugin_rs1Data = 1'b1;
  assign _zz_decode_RegFilePlugin_rs2Data = 1'b1;
  assign _zz_IBusCachedPlugin_jump_pcLoad_payload_6 = {_zz_IBusCachedPlugin_jump_pcLoad_payload_4,_zz_IBusCachedPlugin_jump_pcLoad_payload_3};
  assign _zz_writeBack_DBusCachedPlugin_rspShifted_1 = dataCache_1_io_cpu_writeBack_address[1 : 0];
  assign _zz_writeBack_DBusCachedPlugin_rspShifted_3 = dataCache_1_io_cpu_writeBack_address[1 : 1];
  assign _zz_PmpPlugin_dGuard_hits_0_2 = 4'b0000;
  assign _zz_PmpPlugin_dGuard_hits_0_4 = 4'b0000;
  assign _zz_PmpPlugin_dGuard_hits_1_1 = 4'b0001;
  assign _zz_PmpPlugin_dGuard_hits_1_3 = 4'b0001;
  assign _zz_PmpPlugin_dGuard_hits_2_1 = 4'b0010;
  assign _zz_PmpPlugin_dGuard_hits_2_3 = 4'b0010;
  assign _zz_PmpPlugin_dGuard_hits_3_1 = 4'b0011;
  assign _zz_PmpPlugin_dGuard_hits_3_3 = 4'b0011;
  assign _zz_PmpPlugin_dGuard_hits_4_1 = 4'b0100;
  assign _zz_PmpPlugin_dGuard_hits_4_3 = 4'b0100;
  assign _zz_PmpPlugin_dGuard_hits_5_1 = 4'b0101;
  assign _zz_PmpPlugin_dGuard_hits_5_3 = 4'b0101;
  assign _zz_PmpPlugin_dGuard_hits_6_1 = 4'b0110;
  assign _zz_PmpPlugin_dGuard_hits_6_3 = 4'b0110;
  assign _zz_PmpPlugin_dGuard_hits_7_1 = 4'b0111;
  assign _zz_PmpPlugin_dGuard_hits_7_3 = 4'b0111;
  assign _zz_PmpPlugin_dGuard_hits_8_1 = 4'b1000;
  assign _zz_PmpPlugin_dGuard_hits_8_3 = 4'b1000;
  assign _zz_PmpPlugin_dGuard_hits_9_1 = 4'b1001;
  assign _zz_PmpPlugin_dGuard_hits_9_3 = 4'b1001;
  assign _zz_PmpPlugin_dGuard_hits_10_1 = 4'b1010;
  assign _zz_PmpPlugin_dGuard_hits_10_3 = 4'b1010;
  assign _zz_PmpPlugin_dGuard_hits_11_1 = 4'b1011;
  assign _zz_PmpPlugin_dGuard_hits_11_3 = 4'b1011;
  assign _zz_PmpPlugin_dGuard_hits_12_1 = 4'b1100;
  assign _zz_PmpPlugin_dGuard_hits_12_3 = 4'b1100;
  assign _zz_PmpPlugin_dGuard_hits_13_1 = 4'b1101;
  assign _zz_PmpPlugin_dGuard_hits_13_3 = 4'b1101;
  assign _zz_PmpPlugin_dGuard_hits_14_1 = 4'b1110;
  assign _zz_PmpPlugin_dGuard_hits_14_3 = 4'b1110;
  assign _zz_PmpPlugin_dGuard_hits_15_1 = 4'b1111;
  assign _zz_PmpPlugin_dGuard_hits_15_3 = 4'b1111;
  assign _zz_DBusCachedPlugin_mmuBus_rsp_allowRead_18 = {_zz_DBusCachedPlugin_mmuBus_rsp_allowRead_16,{_zz_DBusCachedPlugin_mmuBus_rsp_allowRead_15,{_zz_DBusCachedPlugin_mmuBus_rsp_allowRead_14,_zz_DBusCachedPlugin_mmuBus_rsp_allowRead_13}}};
  assign _zz_DBusCachedPlugin_mmuBus_rsp_allowWrite_18 = {_zz_DBusCachedPlugin_mmuBus_rsp_allowWrite_16,{_zz_DBusCachedPlugin_mmuBus_rsp_allowWrite_15,{_zz_DBusCachedPlugin_mmuBus_rsp_allowWrite_14,_zz_DBusCachedPlugin_mmuBus_rsp_allowWrite_13}}};
  assign _zz_PmpPlugin_iGuard_hits_0_2 = 4'b0000;
  assign _zz_PmpPlugin_iGuard_hits_0_4 = 4'b0000;
  assign _zz_PmpPlugin_iGuard_hits_1_1 = 4'b0001;
  assign _zz_PmpPlugin_iGuard_hits_1_3 = 4'b0001;
  assign _zz_PmpPlugin_iGuard_hits_2_1 = 4'b0010;
  assign _zz_PmpPlugin_iGuard_hits_2_3 = 4'b0010;
  assign _zz_PmpPlugin_iGuard_hits_3_1 = 4'b0011;
  assign _zz_PmpPlugin_iGuard_hits_3_3 = 4'b0011;
  assign _zz_PmpPlugin_iGuard_hits_4_1 = 4'b0100;
  assign _zz_PmpPlugin_iGuard_hits_4_3 = 4'b0100;
  assign _zz_PmpPlugin_iGuard_hits_5_1 = 4'b0101;
  assign _zz_PmpPlugin_iGuard_hits_5_3 = 4'b0101;
  assign _zz_PmpPlugin_iGuard_hits_6_1 = 4'b0110;
  assign _zz_PmpPlugin_iGuard_hits_6_3 = 4'b0110;
  assign _zz_PmpPlugin_iGuard_hits_7_1 = 4'b0111;
  assign _zz_PmpPlugin_iGuard_hits_7_3 = 4'b0111;
  assign _zz_PmpPlugin_iGuard_hits_8_1 = 4'b1000;
  assign _zz_PmpPlugin_iGuard_hits_8_3 = 4'b1000;
  assign _zz_PmpPlugin_iGuard_hits_9_1 = 4'b1001;
  assign _zz_PmpPlugin_iGuard_hits_9_3 = 4'b1001;
  assign _zz_PmpPlugin_iGuard_hits_10_1 = 4'b1010;
  assign _zz_PmpPlugin_iGuard_hits_10_3 = 4'b1010;
  assign _zz_PmpPlugin_iGuard_hits_11_1 = 4'b1011;
  assign _zz_PmpPlugin_iGuard_hits_11_3 = 4'b1011;
  assign _zz_PmpPlugin_iGuard_hits_12_1 = 4'b1100;
  assign _zz_PmpPlugin_iGuard_hits_12_3 = 4'b1100;
  assign _zz_PmpPlugin_iGuard_hits_13_1 = 4'b1101;
  assign _zz_PmpPlugin_iGuard_hits_13_3 = 4'b1101;
  assign _zz_PmpPlugin_iGuard_hits_14_1 = 4'b1110;
  assign _zz_PmpPlugin_iGuard_hits_14_3 = 4'b1110;
  assign _zz_PmpPlugin_iGuard_hits_15_1 = 4'b1111;
  assign _zz_PmpPlugin_iGuard_hits_15_3 = 4'b1111;
  assign _zz_IBusCachedPlugin_mmuBus_rsp_allowExecute_18 = {_zz_IBusCachedPlugin_mmuBus_rsp_allowExecute_16,{_zz_IBusCachedPlugin_mmuBus_rsp_allowExecute_15,{_zz_IBusCachedPlugin_mmuBus_rsp_allowExecute_14,_zz_IBusCachedPlugin_mmuBus_rsp_allowExecute_13}}};
  assign _zz_when_PmpPlugin_l209_1 = {execute_PmpPlugin_pmpcfgN_,2'b00};
  assign _zz_when_PmpPlugin_l209_1_2 = {execute_PmpPlugin_pmpcfgN_,2'b01};
  assign _zz_when_PmpPlugin_l209_2_1 = {execute_PmpPlugin_pmpcfgN_,2'b10};
  assign _zz_when_PmpPlugin_l209_3_1 = {execute_PmpPlugin_pmpcfgN_,2'b11};
  assign _zz_CsrPlugin_csrMapping_readDataSignal_1 = {execute_PmpPlugin_pmpcfgN,2'b11};
  assign _zz_CsrPlugin_csrMapping_readDataSignal_3 = {execute_PmpPlugin_pmpcfgN,2'b10};
  assign _zz_CsrPlugin_csrMapping_readDataSignal_5 = {execute_PmpPlugin_pmpcfgN,2'b01};
  assign _zz_CsrPlugin_csrMapping_readDataSignal_7 = {execute_PmpPlugin_pmpcfgN,2'b00};
  assign _zz_decode_LEGAL_INSTRUCTION = 32'h0000107f;
  assign _zz_decode_LEGAL_INSTRUCTION_1 = (decode_INSTRUCTION & 32'h0000207f);
  assign _zz_decode_LEGAL_INSTRUCTION_2 = 32'h00002073;
  assign _zz_decode_LEGAL_INSTRUCTION_3 = ((decode_INSTRUCTION & 32'h0000407f) == 32'h00004063);
  assign _zz_decode_LEGAL_INSTRUCTION_4 = ((decode_INSTRUCTION & 32'h0000207f) == 32'h00002013);
  assign _zz_decode_LEGAL_INSTRUCTION_5 = {((decode_INSTRUCTION & 32'h0000603f) == 32'h00000023),{((decode_INSTRUCTION & 32'h0000207f) == 32'h00000003),{((decode_INSTRUCTION & _zz_decode_LEGAL_INSTRUCTION_6) == 32'h00000003),{(_zz_decode_LEGAL_INSTRUCTION_7 == _zz_decode_LEGAL_INSTRUCTION_8),{_zz_decode_LEGAL_INSTRUCTION_9,{_zz_decode_LEGAL_INSTRUCTION_10,_zz_decode_LEGAL_INSTRUCTION_11}}}}}};
  assign _zz_decode_LEGAL_INSTRUCTION_6 = 32'h0000505f;
  assign _zz_decode_LEGAL_INSTRUCTION_7 = (decode_INSTRUCTION & 32'h0000707b);
  assign _zz_decode_LEGAL_INSTRUCTION_8 = 32'h00000063;
  assign _zz_decode_LEGAL_INSTRUCTION_9 = ((decode_INSTRUCTION & 32'h0000607f) == 32'h0000000f);
  assign _zz_decode_LEGAL_INSTRUCTION_10 = ((decode_INSTRUCTION & 32'hfc00007f) == 32'h00000033);
  assign _zz_decode_LEGAL_INSTRUCTION_11 = {((decode_INSTRUCTION & 32'h01f0707f) == 32'h0000500f),{((decode_INSTRUCTION & 32'hbc00707f) == 32'h00005013),{((decode_INSTRUCTION & _zz_decode_LEGAL_INSTRUCTION_12) == 32'h00001013),{(_zz_decode_LEGAL_INSTRUCTION_13 == _zz_decode_LEGAL_INSTRUCTION_14),{_zz_decode_LEGAL_INSTRUCTION_15,{_zz_decode_LEGAL_INSTRUCTION_16,_zz_decode_LEGAL_INSTRUCTION_17}}}}}};
  assign _zz_decode_LEGAL_INSTRUCTION_12 = 32'hfc00307f;
  assign _zz_decode_LEGAL_INSTRUCTION_13 = (decode_INSTRUCTION & 32'hbe00707f);
  assign _zz_decode_LEGAL_INSTRUCTION_14 = 32'h00005033;
  assign _zz_decode_LEGAL_INSTRUCTION_15 = ((decode_INSTRUCTION & 32'hbe00707f) == 32'h00000033);
  assign _zz_decode_LEGAL_INSTRUCTION_16 = ((decode_INSTRUCTION & 32'hdfffffff) == 32'h10200073);
  assign _zz_decode_LEGAL_INSTRUCTION_17 = {((decode_INSTRUCTION & 32'hffffffff) == 32'h10500073),((decode_INSTRUCTION & 32'hffffffff) == 32'h00000073)};
  assign _zz_IBusCachedPlugin_predictionJumpInterface_payload_4 = decode_INSTRUCTION[31];
  assign _zz_IBusCachedPlugin_predictionJumpInterface_payload_5 = decode_INSTRUCTION[31];
  assign _zz_IBusCachedPlugin_predictionJumpInterface_payload_6 = decode_INSTRUCTION[7];
  assign _zz_when_PmpPlugin_l277 = PmpPlugin_dGuard_hits_6;
  assign _zz_when_PmpPlugin_l277_1 = {PmpPlugin_dGuard_hits_5,{PmpPlugin_dGuard_hits_4,{PmpPlugin_dGuard_hits_3,{PmpPlugin_dGuard_hits_2,{PmpPlugin_dGuard_hits_1,PmpPlugin_dGuard_hits_0}}}}};
  assign _zz__zz_DBusCachedPlugin_mmuBus_rsp_allowRead = PmpPlugin_dGuard_hits_5;
  assign _zz__zz_DBusCachedPlugin_mmuBus_rsp_allowRead_1 = {PmpPlugin_dGuard_hits_4,{PmpPlugin_dGuard_hits_3,{PmpPlugin_dGuard_hits_2,{PmpPlugin_dGuard_hits_1,PmpPlugin_dGuard_hits_0}}}};
  assign _zz__zz_DBusCachedPlugin_mmuBus_rsp_allowWrite = PmpPlugin_dGuard_hits_5;
  assign _zz__zz_DBusCachedPlugin_mmuBus_rsp_allowWrite_1 = {PmpPlugin_dGuard_hits_4,{PmpPlugin_dGuard_hits_3,{PmpPlugin_dGuard_hits_2,{PmpPlugin_dGuard_hits_1,PmpPlugin_dGuard_hits_0}}}};
  assign _zz_when_PmpPlugin_l299 = PmpPlugin_iGuard_hits_6;
  assign _zz_when_PmpPlugin_l299_1 = {PmpPlugin_iGuard_hits_5,{PmpPlugin_iGuard_hits_4,{PmpPlugin_iGuard_hits_3,{PmpPlugin_iGuard_hits_2,{PmpPlugin_iGuard_hits_1,PmpPlugin_iGuard_hits_0}}}}};
  assign _zz__zz_IBusCachedPlugin_mmuBus_rsp_allowExecute = PmpPlugin_iGuard_hits_5;
  assign _zz__zz_IBusCachedPlugin_mmuBus_rsp_allowExecute_1 = {PmpPlugin_iGuard_hits_4,{PmpPlugin_iGuard_hits_3,{PmpPlugin_iGuard_hits_2,{PmpPlugin_iGuard_hits_1,PmpPlugin_iGuard_hits_0}}}};
  assign _zz__zz_decode_IS_RS2_SIGNED = (decode_INSTRUCTION & 32'h02004064);
  assign _zz__zz_decode_IS_RS2_SIGNED_1 = 32'h02004020;
  assign _zz__zz_decode_IS_RS2_SIGNED_2 = ((decode_INSTRUCTION & 32'h02004074) == 32'h02000030);
  assign _zz__zz_decode_IS_RS2_SIGNED_3 = ((decode_INSTRUCTION & 32'h00203050) == 32'h00000050);
  assign _zz__zz_decode_IS_RS2_SIGNED_4 = (|((decode_INSTRUCTION & _zz__zz_decode_IS_RS2_SIGNED_5) == 32'h00000050));
  assign _zz__zz_decode_IS_RS2_SIGNED_6 = (|{_zz__zz_decode_IS_RS2_SIGNED_7,_zz__zz_decode_IS_RS2_SIGNED_8});
  assign _zz__zz_decode_IS_RS2_SIGNED_9 = {(|{_zz__zz_decode_IS_RS2_SIGNED_10,_zz__zz_decode_IS_RS2_SIGNED_11}),{(|_zz__zz_decode_IS_RS2_SIGNED_13),{_zz__zz_decode_IS_RS2_SIGNED_15,{_zz__zz_decode_IS_RS2_SIGNED_18,_zz__zz_decode_IS_RS2_SIGNED_26}}}};
  assign _zz__zz_decode_IS_RS2_SIGNED_5 = 32'h00403050;
  assign _zz__zz_decode_IS_RS2_SIGNED_7 = ((decode_INSTRUCTION & 32'h00001050) == 32'h00001050);
  assign _zz__zz_decode_IS_RS2_SIGNED_8 = ((decode_INSTRUCTION & 32'h00002050) == 32'h00002050);
  assign _zz__zz_decode_IS_RS2_SIGNED_10 = _zz_decode_IS_RS2_SIGNED_4;
  assign _zz__zz_decode_IS_RS2_SIGNED_11 = ((decode_INSTRUCTION & _zz__zz_decode_IS_RS2_SIGNED_12) == 32'h00000004);
  assign _zz__zz_decode_IS_RS2_SIGNED_13 = ((decode_INSTRUCTION & _zz__zz_decode_IS_RS2_SIGNED_14) == 32'h00000040);
  assign _zz__zz_decode_IS_RS2_SIGNED_15 = (|{_zz__zz_decode_IS_RS2_SIGNED_16,_zz__zz_decode_IS_RS2_SIGNED_17});
  assign _zz__zz_decode_IS_RS2_SIGNED_18 = (|{_zz__zz_decode_IS_RS2_SIGNED_19,_zz__zz_decode_IS_RS2_SIGNED_21});
  assign _zz__zz_decode_IS_RS2_SIGNED_26 = {(|_zz__zz_decode_IS_RS2_SIGNED_27),{_zz__zz_decode_IS_RS2_SIGNED_29,{_zz__zz_decode_IS_RS2_SIGNED_32,_zz__zz_decode_IS_RS2_SIGNED_34}}};
  assign _zz__zz_decode_IS_RS2_SIGNED_12 = 32'h0000001c;
  assign _zz__zz_decode_IS_RS2_SIGNED_14 = 32'h00000058;
  assign _zz__zz_decode_IS_RS2_SIGNED_16 = ((decode_INSTRUCTION & 32'h00007034) == 32'h00005010);
  assign _zz__zz_decode_IS_RS2_SIGNED_17 = ((decode_INSTRUCTION & 32'h02007064) == 32'h00005020);
  assign _zz__zz_decode_IS_RS2_SIGNED_19 = ((decode_INSTRUCTION & _zz__zz_decode_IS_RS2_SIGNED_20) == 32'h40001010);
  assign _zz__zz_decode_IS_RS2_SIGNED_21 = {(_zz__zz_decode_IS_RS2_SIGNED_22 == _zz__zz_decode_IS_RS2_SIGNED_23),(_zz__zz_decode_IS_RS2_SIGNED_24 == _zz__zz_decode_IS_RS2_SIGNED_25)};
  assign _zz__zz_decode_IS_RS2_SIGNED_27 = ((decode_INSTRUCTION & _zz__zz_decode_IS_RS2_SIGNED_28) == 32'h00000024);
  assign _zz__zz_decode_IS_RS2_SIGNED_29 = (|(_zz__zz_decode_IS_RS2_SIGNED_30 == _zz__zz_decode_IS_RS2_SIGNED_31));
  assign _zz__zz_decode_IS_RS2_SIGNED_32 = (|_zz__zz_decode_IS_RS2_SIGNED_33);
  assign _zz__zz_decode_IS_RS2_SIGNED_34 = {(|_zz__zz_decode_IS_RS2_SIGNED_35),{_zz__zz_decode_IS_RS2_SIGNED_38,{_zz__zz_decode_IS_RS2_SIGNED_40,_zz__zz_decode_IS_RS2_SIGNED_43}}};
  assign _zz__zz_decode_IS_RS2_SIGNED_20 = 32'h40003054;
  assign _zz__zz_decode_IS_RS2_SIGNED_22 = (decode_INSTRUCTION & 32'h00007034);
  assign _zz__zz_decode_IS_RS2_SIGNED_23 = 32'h00001010;
  assign _zz__zz_decode_IS_RS2_SIGNED_24 = (decode_INSTRUCTION & 32'h02007054);
  assign _zz__zz_decode_IS_RS2_SIGNED_25 = 32'h00001010;
  assign _zz__zz_decode_IS_RS2_SIGNED_28 = 32'h00000064;
  assign _zz__zz_decode_IS_RS2_SIGNED_30 = (decode_INSTRUCTION & 32'h00001000);
  assign _zz__zz_decode_IS_RS2_SIGNED_31 = 32'h00001000;
  assign _zz__zz_decode_IS_RS2_SIGNED_33 = ((decode_INSTRUCTION & 32'h00003000) == 32'h00002000);
  assign _zz__zz_decode_IS_RS2_SIGNED_35 = {((decode_INSTRUCTION & _zz__zz_decode_IS_RS2_SIGNED_36) == 32'h00002000),((decode_INSTRUCTION & _zz__zz_decode_IS_RS2_SIGNED_37) == 32'h00001000)};
  assign _zz__zz_decode_IS_RS2_SIGNED_38 = (|((decode_INSTRUCTION & _zz__zz_decode_IS_RS2_SIGNED_39) == 32'h00004008));
  assign _zz__zz_decode_IS_RS2_SIGNED_40 = (|{_zz__zz_decode_IS_RS2_SIGNED_41,_zz__zz_decode_IS_RS2_SIGNED_42});
  assign _zz__zz_decode_IS_RS2_SIGNED_43 = {(|{_zz__zz_decode_IS_RS2_SIGNED_44,_zz__zz_decode_IS_RS2_SIGNED_46}),{(|_zz__zz_decode_IS_RS2_SIGNED_55),{_zz__zz_decode_IS_RS2_SIGNED_57,{_zz__zz_decode_IS_RS2_SIGNED_70,_zz__zz_decode_IS_RS2_SIGNED_83}}}};
  assign _zz__zz_decode_IS_RS2_SIGNED_36 = 32'h00002010;
  assign _zz__zz_decode_IS_RS2_SIGNED_37 = 32'h00005000;
  assign _zz__zz_decode_IS_RS2_SIGNED_39 = 32'h00004048;
  assign _zz__zz_decode_IS_RS2_SIGNED_41 = ((decode_INSTRUCTION & 32'h00000034) == 32'h00000020);
  assign _zz__zz_decode_IS_RS2_SIGNED_42 = ((decode_INSTRUCTION & 32'h00000064) == 32'h00000020);
  assign _zz__zz_decode_IS_RS2_SIGNED_44 = ((decode_INSTRUCTION & _zz__zz_decode_IS_RS2_SIGNED_45) == 32'h00002040);
  assign _zz__zz_decode_IS_RS2_SIGNED_46 = {(_zz__zz_decode_IS_RS2_SIGNED_47 == _zz__zz_decode_IS_RS2_SIGNED_48),{_zz__zz_decode_IS_RS2_SIGNED_49,{_zz__zz_decode_IS_RS2_SIGNED_51,_zz__zz_decode_IS_RS2_SIGNED_54}}};
  assign _zz__zz_decode_IS_RS2_SIGNED_55 = ((decode_INSTRUCTION & _zz__zz_decode_IS_RS2_SIGNED_56) == 32'h00000020);
  assign _zz__zz_decode_IS_RS2_SIGNED_57 = (|{_zz__zz_decode_IS_RS2_SIGNED_58,{_zz__zz_decode_IS_RS2_SIGNED_60,_zz__zz_decode_IS_RS2_SIGNED_61}});
  assign _zz__zz_decode_IS_RS2_SIGNED_70 = (|{_zz__zz_decode_IS_RS2_SIGNED_71,_zz__zz_decode_IS_RS2_SIGNED_72});
  assign _zz__zz_decode_IS_RS2_SIGNED_83 = {(|_zz__zz_decode_IS_RS2_SIGNED_84),{_zz__zz_decode_IS_RS2_SIGNED_97,{_zz__zz_decode_IS_RS2_SIGNED_102,_zz__zz_decode_IS_RS2_SIGNED_106}}};
  assign _zz__zz_decode_IS_RS2_SIGNED_45 = 32'h00002040;
  assign _zz__zz_decode_IS_RS2_SIGNED_47 = (decode_INSTRUCTION & 32'h00001040);
  assign _zz__zz_decode_IS_RS2_SIGNED_48 = 32'h00001040;
  assign _zz__zz_decode_IS_RS2_SIGNED_49 = ((decode_INSTRUCTION & _zz__zz_decode_IS_RS2_SIGNED_50) == 32'h00000040);
  assign _zz__zz_decode_IS_RS2_SIGNED_51 = (_zz__zz_decode_IS_RS2_SIGNED_52 == _zz__zz_decode_IS_RS2_SIGNED_53);
  assign _zz__zz_decode_IS_RS2_SIGNED_54 = _zz_decode_IS_RS2_SIGNED_2;
  assign _zz__zz_decode_IS_RS2_SIGNED_56 = 32'h00000020;
  assign _zz__zz_decode_IS_RS2_SIGNED_58 = ((decode_INSTRUCTION & _zz__zz_decode_IS_RS2_SIGNED_59) == 32'h00000040);
  assign _zz__zz_decode_IS_RS2_SIGNED_60 = _zz_decode_IS_RS2_SIGNED_3;
  assign _zz__zz_decode_IS_RS2_SIGNED_61 = {_zz__zz_decode_IS_RS2_SIGNED_62,{_zz__zz_decode_IS_RS2_SIGNED_64,_zz__zz_decode_IS_RS2_SIGNED_67}};
  assign _zz__zz_decode_IS_RS2_SIGNED_71 = _zz_decode_IS_RS2_SIGNED_3;
  assign _zz__zz_decode_IS_RS2_SIGNED_72 = {_zz__zz_decode_IS_RS2_SIGNED_73,{_zz__zz_decode_IS_RS2_SIGNED_75,_zz__zz_decode_IS_RS2_SIGNED_78}};
  assign _zz__zz_decode_IS_RS2_SIGNED_84 = {_zz_decode_IS_RS2_SIGNED_4,{_zz__zz_decode_IS_RS2_SIGNED_85,_zz__zz_decode_IS_RS2_SIGNED_88}};
  assign _zz__zz_decode_IS_RS2_SIGNED_97 = (|{_zz__zz_decode_IS_RS2_SIGNED_98,_zz__zz_decode_IS_RS2_SIGNED_99});
  assign _zz__zz_decode_IS_RS2_SIGNED_102 = (|_zz__zz_decode_IS_RS2_SIGNED_103);
  assign _zz__zz_decode_IS_RS2_SIGNED_106 = {_zz__zz_decode_IS_RS2_SIGNED_107,{_zz__zz_decode_IS_RS2_SIGNED_110,_zz__zz_decode_IS_RS2_SIGNED_114}};
  assign _zz__zz_decode_IS_RS2_SIGNED_50 = 32'h00000050;
  assign _zz__zz_decode_IS_RS2_SIGNED_52 = (decode_INSTRUCTION & 32'h00400040);
  assign _zz__zz_decode_IS_RS2_SIGNED_53 = 32'h00000040;
  assign _zz__zz_decode_IS_RS2_SIGNED_59 = 32'h00000040;
  assign _zz__zz_decode_IS_RS2_SIGNED_62 = ((decode_INSTRUCTION & _zz__zz_decode_IS_RS2_SIGNED_63) == 32'h00004020);
  assign _zz__zz_decode_IS_RS2_SIGNED_64 = (_zz__zz_decode_IS_RS2_SIGNED_65 == _zz__zz_decode_IS_RS2_SIGNED_66);
  assign _zz__zz_decode_IS_RS2_SIGNED_67 = (_zz__zz_decode_IS_RS2_SIGNED_68 == _zz__zz_decode_IS_RS2_SIGNED_69);
  assign _zz__zz_decode_IS_RS2_SIGNED_73 = ((decode_INSTRUCTION & _zz__zz_decode_IS_RS2_SIGNED_74) == 32'h00002010);
  assign _zz__zz_decode_IS_RS2_SIGNED_75 = (_zz__zz_decode_IS_RS2_SIGNED_76 == _zz__zz_decode_IS_RS2_SIGNED_77);
  assign _zz__zz_decode_IS_RS2_SIGNED_78 = {_zz__zz_decode_IS_RS2_SIGNED_79,_zz__zz_decode_IS_RS2_SIGNED_81};
  assign _zz__zz_decode_IS_RS2_SIGNED_85 = (_zz__zz_decode_IS_RS2_SIGNED_86 == _zz__zz_decode_IS_RS2_SIGNED_87);
  assign _zz__zz_decode_IS_RS2_SIGNED_88 = {_zz__zz_decode_IS_RS2_SIGNED_89,{_zz__zz_decode_IS_RS2_SIGNED_91,_zz__zz_decode_IS_RS2_SIGNED_94}};
  assign _zz__zz_decode_IS_RS2_SIGNED_98 = _zz_decode_IS_RS2_SIGNED_3;
  assign _zz__zz_decode_IS_RS2_SIGNED_99 = (_zz__zz_decode_IS_RS2_SIGNED_100 == _zz__zz_decode_IS_RS2_SIGNED_101);
  assign _zz__zz_decode_IS_RS2_SIGNED_103 = {_zz_decode_IS_RS2_SIGNED_3,_zz__zz_decode_IS_RS2_SIGNED_104};
  assign _zz__zz_decode_IS_RS2_SIGNED_107 = (|_zz__zz_decode_IS_RS2_SIGNED_108);
  assign _zz__zz_decode_IS_RS2_SIGNED_110 = (|_zz__zz_decode_IS_RS2_SIGNED_111);
  assign _zz__zz_decode_IS_RS2_SIGNED_114 = {_zz__zz_decode_IS_RS2_SIGNED_115,{_zz__zz_decode_IS_RS2_SIGNED_124,_zz__zz_decode_IS_RS2_SIGNED_127}};
  assign _zz__zz_decode_IS_RS2_SIGNED_63 = 32'h00004020;
  assign _zz__zz_decode_IS_RS2_SIGNED_65 = (decode_INSTRUCTION & 32'h00000030);
  assign _zz__zz_decode_IS_RS2_SIGNED_66 = 32'h00000010;
  assign _zz__zz_decode_IS_RS2_SIGNED_68 = (decode_INSTRUCTION & 32'h02000020);
  assign _zz__zz_decode_IS_RS2_SIGNED_69 = 32'h00000020;
  assign _zz__zz_decode_IS_RS2_SIGNED_74 = 32'h00002030;
  assign _zz__zz_decode_IS_RS2_SIGNED_76 = (decode_INSTRUCTION & 32'h00001030);
  assign _zz__zz_decode_IS_RS2_SIGNED_77 = 32'h00000010;
  assign _zz__zz_decode_IS_RS2_SIGNED_79 = ((decode_INSTRUCTION & _zz__zz_decode_IS_RS2_SIGNED_80) == 32'h00002020);
  assign _zz__zz_decode_IS_RS2_SIGNED_81 = ((decode_INSTRUCTION & _zz__zz_decode_IS_RS2_SIGNED_82) == 32'h00000020);
  assign _zz__zz_decode_IS_RS2_SIGNED_86 = (decode_INSTRUCTION & 32'h00001010);
  assign _zz__zz_decode_IS_RS2_SIGNED_87 = 32'h00001010;
  assign _zz__zz_decode_IS_RS2_SIGNED_89 = ((decode_INSTRUCTION & _zz__zz_decode_IS_RS2_SIGNED_90) == 32'h00002010);
  assign _zz__zz_decode_IS_RS2_SIGNED_91 = (_zz__zz_decode_IS_RS2_SIGNED_92 == _zz__zz_decode_IS_RS2_SIGNED_93);
  assign _zz__zz_decode_IS_RS2_SIGNED_94 = {_zz__zz_decode_IS_RS2_SIGNED_95,_zz__zz_decode_IS_RS2_SIGNED_96};
  assign _zz__zz_decode_IS_RS2_SIGNED_100 = (decode_INSTRUCTION & 32'h00000070);
  assign _zz__zz_decode_IS_RS2_SIGNED_101 = 32'h00000020;
  assign _zz__zz_decode_IS_RS2_SIGNED_104 = ((decode_INSTRUCTION & _zz__zz_decode_IS_RS2_SIGNED_105) == 32'h0);
  assign _zz__zz_decode_IS_RS2_SIGNED_108 = ((decode_INSTRUCTION & _zz__zz_decode_IS_RS2_SIGNED_109) == 32'h00004010);
  assign _zz__zz_decode_IS_RS2_SIGNED_111 = (_zz__zz_decode_IS_RS2_SIGNED_112 == _zz__zz_decode_IS_RS2_SIGNED_113);
  assign _zz__zz_decode_IS_RS2_SIGNED_115 = (|{_zz__zz_decode_IS_RS2_SIGNED_116,_zz__zz_decode_IS_RS2_SIGNED_118});
  assign _zz__zz_decode_IS_RS2_SIGNED_124 = (|_zz__zz_decode_IS_RS2_SIGNED_125);
  assign _zz__zz_decode_IS_RS2_SIGNED_127 = {_zz__zz_decode_IS_RS2_SIGNED_128,{_zz__zz_decode_IS_RS2_SIGNED_134,_zz__zz_decode_IS_RS2_SIGNED_138}};
  assign _zz__zz_decode_IS_RS2_SIGNED_80 = 32'h02002060;
  assign _zz__zz_decode_IS_RS2_SIGNED_82 = 32'h02003020;
  assign _zz__zz_decode_IS_RS2_SIGNED_90 = 32'h00002010;
  assign _zz__zz_decode_IS_RS2_SIGNED_92 = (decode_INSTRUCTION & 32'h00000050);
  assign _zz__zz_decode_IS_RS2_SIGNED_93 = 32'h00000010;
  assign _zz__zz_decode_IS_RS2_SIGNED_95 = ((decode_INSTRUCTION & 32'h0000000c) == 32'h00000004);
  assign _zz__zz_decode_IS_RS2_SIGNED_96 = ((decode_INSTRUCTION & 32'h00000028) == 32'h0);
  assign _zz__zz_decode_IS_RS2_SIGNED_105 = 32'h00000020;
  assign _zz__zz_decode_IS_RS2_SIGNED_109 = 32'h00004014;
  assign _zz__zz_decode_IS_RS2_SIGNED_112 = (decode_INSTRUCTION & 32'h00006014);
  assign _zz__zz_decode_IS_RS2_SIGNED_113 = 32'h00002010;
  assign _zz__zz_decode_IS_RS2_SIGNED_116 = ((decode_INSTRUCTION & _zz__zz_decode_IS_RS2_SIGNED_117) == 32'h0);
  assign _zz__zz_decode_IS_RS2_SIGNED_118 = {_zz_decode_IS_RS2_SIGNED_2,{_zz__zz_decode_IS_RS2_SIGNED_119,{_zz__zz_decode_IS_RS2_SIGNED_120,_zz__zz_decode_IS_RS2_SIGNED_122}}};
  assign _zz__zz_decode_IS_RS2_SIGNED_125 = ((decode_INSTRUCTION & _zz__zz_decode_IS_RS2_SIGNED_126) == 32'h0);
  assign _zz__zz_decode_IS_RS2_SIGNED_128 = (|{_zz__zz_decode_IS_RS2_SIGNED_129,{_zz__zz_decode_IS_RS2_SIGNED_130,_zz__zz_decode_IS_RS2_SIGNED_132}});
  assign _zz__zz_decode_IS_RS2_SIGNED_134 = (|{_zz__zz_decode_IS_RS2_SIGNED_135,_zz__zz_decode_IS_RS2_SIGNED_137});
  assign _zz__zz_decode_IS_RS2_SIGNED_138 = {(|_zz__zz_decode_IS_RS2_SIGNED_139),(|_zz__zz_decode_IS_RS2_SIGNED_142)};
  assign _zz__zz_decode_IS_RS2_SIGNED_117 = 32'h00000044;
  assign _zz__zz_decode_IS_RS2_SIGNED_119 = ((decode_INSTRUCTION & 32'h00006004) == 32'h00002000);
  assign _zz__zz_decode_IS_RS2_SIGNED_120 = ((decode_INSTRUCTION & _zz__zz_decode_IS_RS2_SIGNED_121) == 32'h00001000);
  assign _zz__zz_decode_IS_RS2_SIGNED_122 = ((decode_INSTRUCTION & _zz__zz_decode_IS_RS2_SIGNED_123) == 32'h00004000);
  assign _zz__zz_decode_IS_RS2_SIGNED_126 = 32'h00000058;
  assign _zz__zz_decode_IS_RS2_SIGNED_129 = ((decode_INSTRUCTION & 32'h00000044) == 32'h00000040);
  assign _zz__zz_decode_IS_RS2_SIGNED_130 = ((decode_INSTRUCTION & _zz__zz_decode_IS_RS2_SIGNED_131) == 32'h00002010);
  assign _zz__zz_decode_IS_RS2_SIGNED_132 = ((decode_INSTRUCTION & _zz__zz_decode_IS_RS2_SIGNED_133) == 32'h40000030);
  assign _zz__zz_decode_IS_RS2_SIGNED_135 = ((decode_INSTRUCTION & _zz__zz_decode_IS_RS2_SIGNED_136) == 32'h00000004);
  assign _zz__zz_decode_IS_RS2_SIGNED_137 = _zz_decode_IS_RS2_SIGNED_1;
  assign _zz__zz_decode_IS_RS2_SIGNED_139 = {(_zz__zz_decode_IS_RS2_SIGNED_140 == _zz__zz_decode_IS_RS2_SIGNED_141),_zz_decode_IS_RS2_SIGNED_1};
  assign _zz__zz_decode_IS_RS2_SIGNED_142 = ((decode_INSTRUCTION & _zz__zz_decode_IS_RS2_SIGNED_143) == 32'h00001008);
  assign _zz__zz_decode_IS_RS2_SIGNED_121 = 32'h00005004;
  assign _zz__zz_decode_IS_RS2_SIGNED_123 = 32'h00004050;
  assign _zz__zz_decode_IS_RS2_SIGNED_131 = 32'h00002014;
  assign _zz__zz_decode_IS_RS2_SIGNED_133 = 32'h40000034;
  assign _zz__zz_decode_IS_RS2_SIGNED_136 = 32'h00000014;
  assign _zz__zz_decode_IS_RS2_SIGNED_140 = (decode_INSTRUCTION & 32'h00000044);
  assign _zz__zz_decode_IS_RS2_SIGNED_141 = 32'h00000004;
  assign _zz__zz_decode_IS_RS2_SIGNED_143 = 32'h00005048;
  assign _zz_execute_BranchPlugin_branch_src2_6 = execute_INSTRUCTION[31];
  assign _zz_execute_BranchPlugin_branch_src2_7 = execute_INSTRUCTION[31];
  assign _zz_execute_BranchPlugin_branch_src2_8 = execute_INSTRUCTION[7];
  assign _zz_CsrPlugin_csrMapping_readDataInit_25 = 32'h0;
  assign _zz_PmpPlugin_pmpaddr_port0 = PmpPlugin_pmpaddr[execute_PmpPlugin_fsm_fsmCounter];
  always @(posedge clk) begin
    if(_zz_1) begin
      PmpPlugin_pmpaddr[execute_PmpPlugin_pmpNcfg_] <= _zz_PmpPlugin_pmpaddr_port;
    end
  end

  assign _zz_PmpPlugin_pmpaddr_port2 = PmpPlugin_pmpaddr[execute_PmpPlugin_pmpNcfg];
  always @(posedge clk) begin
    if(_zz_decode_RegFilePlugin_rs1Data) begin
      _zz_RegFilePlugin_regFile_port0 <= RegFilePlugin_regFile[decode_RegFilePlugin_regFileReadAddress1];
    end
  end

  always @(posedge clk) begin
    if(_zz_decode_RegFilePlugin_rs2Data) begin
      _zz_RegFilePlugin_regFile_port1 <= RegFilePlugin_regFile[decode_RegFilePlugin_regFileReadAddress2];
    end
  end

  always @(posedge clk) begin
    if(_zz_2) begin
      RegFilePlugin_regFile[lastStageRegFileWrite_payload_address] <= lastStageRegFileWrite_payload_data;
    end
  end

  PmpSetter PmpPlugin_setter (
    .io_addr (PmpPlugin_setter_io_addr[31:0]), //i
    .io_base (PmpPlugin_setter_io_base[24:0]), //o
    .io_mask (PmpPlugin_setter_io_mask[24:0])  //o
  );
  InstructionCache IBusCachedPlugin_cache (
    .io_flush                              (IBusCachedPlugin_cache_io_flush                           ), //i
    .io_cpu_prefetch_isValid               (IBusCachedPlugin_cache_io_cpu_prefetch_isValid            ), //i
    .io_cpu_prefetch_haltIt                (IBusCachedPlugin_cache_io_cpu_prefetch_haltIt             ), //o
    .io_cpu_prefetch_pc                    (IBusCachedPlugin_iBusRsp_stages_0_input_payload[31:0]     ), //i
    .io_cpu_fetch_isValid                  (IBusCachedPlugin_cache_io_cpu_fetch_isValid               ), //i
    .io_cpu_fetch_isStuck                  (IBusCachedPlugin_cache_io_cpu_fetch_isStuck               ), //i
    .io_cpu_fetch_isRemoved                (IBusCachedPlugin_cache_io_cpu_fetch_isRemoved             ), //i
    .io_cpu_fetch_pc                       (IBusCachedPlugin_iBusRsp_stages_1_input_payload[31:0]     ), //i
    .io_cpu_fetch_data                     (IBusCachedPlugin_cache_io_cpu_fetch_data[31:0]            ), //o
    .io_cpu_fetch_mmuRsp_physicalAddress   (IBusCachedPlugin_mmuBus_rsp_physicalAddress[31:0]         ), //i
    .io_cpu_fetch_mmuRsp_isIoAccess        (IBusCachedPlugin_mmuBus_rsp_isIoAccess                    ), //i
    .io_cpu_fetch_mmuRsp_isPaging          (IBusCachedPlugin_mmuBus_rsp_isPaging                      ), //i
    .io_cpu_fetch_mmuRsp_allowRead         (IBusCachedPlugin_mmuBus_rsp_allowRead                     ), //i
    .io_cpu_fetch_mmuRsp_allowWrite        (IBusCachedPlugin_mmuBus_rsp_allowWrite                    ), //i
    .io_cpu_fetch_mmuRsp_allowExecute      (IBusCachedPlugin_mmuBus_rsp_allowExecute                  ), //i
    .io_cpu_fetch_mmuRsp_exception         (IBusCachedPlugin_mmuBus_rsp_exception                     ), //i
    .io_cpu_fetch_mmuRsp_refilling         (IBusCachedPlugin_mmuBus_rsp_refilling                     ), //i
    .io_cpu_fetch_mmuRsp_bypassTranslation (IBusCachedPlugin_mmuBus_rsp_bypassTranslation             ), //i
    .io_cpu_fetch_physicalAddress          (IBusCachedPlugin_cache_io_cpu_fetch_physicalAddress[31:0] ), //o
    .io_cpu_decode_isValid                 (IBusCachedPlugin_cache_io_cpu_decode_isValid              ), //i
    .io_cpu_decode_isStuck                 (IBusCachedPlugin_cache_io_cpu_decode_isStuck              ), //i
    .io_cpu_decode_pc                      (IBusCachedPlugin_iBusRsp_stages_2_input_payload[31:0]     ), //i
    .io_cpu_decode_physicalAddress         (IBusCachedPlugin_cache_io_cpu_decode_physicalAddress[31:0]), //o
    .io_cpu_decode_data                    (IBusCachedPlugin_cache_io_cpu_decode_data[31:0]           ), //o
    .io_cpu_decode_cacheMiss               (IBusCachedPlugin_cache_io_cpu_decode_cacheMiss            ), //o
    .io_cpu_decode_error                   (IBusCachedPlugin_cache_io_cpu_decode_error                ), //o
    .io_cpu_decode_mmuRefilling            (IBusCachedPlugin_cache_io_cpu_decode_mmuRefilling         ), //o
    .io_cpu_decode_mmuException            (IBusCachedPlugin_cache_io_cpu_decode_mmuException         ), //o
    .io_cpu_decode_isUser                  (IBusCachedPlugin_cache_io_cpu_decode_isUser               ), //i
    .io_cpu_fill_valid                     (IBusCachedPlugin_cache_io_cpu_fill_valid                  ), //i
    .io_cpu_fill_payload                   (IBusCachedPlugin_cache_io_cpu_decode_physicalAddress[31:0]), //i
    .io_mem_cmd_valid                      (IBusCachedPlugin_cache_io_mem_cmd_valid                   ), //o
    .io_mem_cmd_ready                      (iBus_cmd_ready                                            ), //i
    .io_mem_cmd_payload_address            (IBusCachedPlugin_cache_io_mem_cmd_payload_address[31:0]   ), //o
    .io_mem_cmd_payload_size               (IBusCachedPlugin_cache_io_mem_cmd_payload_size[2:0]       ), //o
    .io_mem_rsp_valid                      (iBus_rsp_valid                                            ), //i
    .io_mem_rsp_payload_data               (iBus_rsp_payload_data[31:0]                               ), //i
    .io_mem_rsp_payload_error              (iBus_rsp_payload_error                                    ), //i
    .clk                                   (clk                                                       ), //i
    .reset                                 (reset                                                     )  //i
  );
  DataCache dataCache_1 (
    .io_cpu_execute_isValid                 (dataCache_1_io_cpu_execute_isValid               ), //i
    .io_cpu_execute_address                 (dataCache_1_io_cpu_execute_address[31:0]         ), //i
    .io_cpu_execute_haltIt                  (dataCache_1_io_cpu_execute_haltIt                ), //o
    .io_cpu_execute_args_wr                 (execute_MEMORY_WR                                ), //i
    .io_cpu_execute_args_size               (execute_DBusCachedPlugin_size[1:0]               ), //i
    .io_cpu_execute_args_totalyConsistent   (execute_MEMORY_FORCE_CONSTISTENCY                ), //i
    .io_cpu_execute_refilling               (dataCache_1_io_cpu_execute_refilling             ), //o
    .io_cpu_memory_isValid                  (dataCache_1_io_cpu_memory_isValid                ), //i
    .io_cpu_memory_isStuck                  (memory_arbitration_isStuck                       ), //i
    .io_cpu_memory_isWrite                  (dataCache_1_io_cpu_memory_isWrite                ), //o
    .io_cpu_memory_address                  (dataCache_1_io_cpu_memory_address[31:0]          ), //i
    .io_cpu_memory_mmuRsp_physicalAddress   (DBusCachedPlugin_mmuBus_rsp_physicalAddress[31:0]), //i
    .io_cpu_memory_mmuRsp_isIoAccess        (dataCache_1_io_cpu_memory_mmuRsp_isIoAccess      ), //i
    .io_cpu_memory_mmuRsp_isPaging          (DBusCachedPlugin_mmuBus_rsp_isPaging             ), //i
    .io_cpu_memory_mmuRsp_allowRead         (DBusCachedPlugin_mmuBus_rsp_allowRead            ), //i
    .io_cpu_memory_mmuRsp_allowWrite        (DBusCachedPlugin_mmuBus_rsp_allowWrite           ), //i
    .io_cpu_memory_mmuRsp_allowExecute      (DBusCachedPlugin_mmuBus_rsp_allowExecute         ), //i
    .io_cpu_memory_mmuRsp_exception         (DBusCachedPlugin_mmuBus_rsp_exception            ), //i
    .io_cpu_memory_mmuRsp_refilling         (DBusCachedPlugin_mmuBus_rsp_refilling            ), //i
    .io_cpu_memory_mmuRsp_bypassTranslation (DBusCachedPlugin_mmuBus_rsp_bypassTranslation    ), //i
    .io_cpu_writeBack_isValid               (dataCache_1_io_cpu_writeBack_isValid             ), //i
    .io_cpu_writeBack_isStuck               (writeBack_arbitration_isStuck                    ), //i
    .io_cpu_writeBack_isFiring              (writeBack_arbitration_isFiring                   ), //i
    .io_cpu_writeBack_isUser                (dataCache_1_io_cpu_writeBack_isUser              ), //i
    .io_cpu_writeBack_haltIt                (dataCache_1_io_cpu_writeBack_haltIt              ), //o
    .io_cpu_writeBack_isWrite               (dataCache_1_io_cpu_writeBack_isWrite             ), //o
    .io_cpu_writeBack_storeData             (dataCache_1_io_cpu_writeBack_storeData[31:0]     ), //i
    .io_cpu_writeBack_data                  (dataCache_1_io_cpu_writeBack_data[31:0]          ), //o
    .io_cpu_writeBack_address               (dataCache_1_io_cpu_writeBack_address[31:0]       ), //i
    .io_cpu_writeBack_mmuException          (dataCache_1_io_cpu_writeBack_mmuException        ), //o
    .io_cpu_writeBack_unalignedAccess       (dataCache_1_io_cpu_writeBack_unalignedAccess     ), //o
    .io_cpu_writeBack_accessError           (dataCache_1_io_cpu_writeBack_accessError         ), //o
    .io_cpu_writeBack_keepMemRspData        (dataCache_1_io_cpu_writeBack_keepMemRspData      ), //o
    .io_cpu_writeBack_fence_SW              (dataCache_1_io_cpu_writeBack_fence_SW            ), //i
    .io_cpu_writeBack_fence_SR              (dataCache_1_io_cpu_writeBack_fence_SR            ), //i
    .io_cpu_writeBack_fence_SO              (dataCache_1_io_cpu_writeBack_fence_SO            ), //i
    .io_cpu_writeBack_fence_SI              (dataCache_1_io_cpu_writeBack_fence_SI            ), //i
    .io_cpu_writeBack_fence_PW              (dataCache_1_io_cpu_writeBack_fence_PW            ), //i
    .io_cpu_writeBack_fence_PR              (dataCache_1_io_cpu_writeBack_fence_PR            ), //i
    .io_cpu_writeBack_fence_PO              (dataCache_1_io_cpu_writeBack_fence_PO            ), //i
    .io_cpu_writeBack_fence_PI              (dataCache_1_io_cpu_writeBack_fence_PI            ), //i
    .io_cpu_writeBack_fence_FM              (dataCache_1_io_cpu_writeBack_fence_FM[3:0]       ), //i
    .io_cpu_writeBack_exclusiveOk           (dataCache_1_io_cpu_writeBack_exclusiveOk         ), //o
    .io_cpu_redo                            (dataCache_1_io_cpu_redo                          ), //o
    .io_cpu_flush_valid                     (dataCache_1_io_cpu_flush_valid                   ), //i
    .io_cpu_flush_ready                     (dataCache_1_io_cpu_flush_ready                   ), //o
    .io_cpu_flush_payload_singleLine        (dataCache_1_io_cpu_flush_payload_singleLine      ), //i
    .io_cpu_flush_payload_lineId            (dataCache_1_io_cpu_flush_payload_lineId[6:0]     ), //i
    .io_mem_cmd_valid                       (dataCache_1_io_mem_cmd_valid                     ), //o
    .io_mem_cmd_ready                       (dataCache_1_io_mem_cmd_ready                     ), //i
    .io_mem_cmd_payload_wr                  (dataCache_1_io_mem_cmd_payload_wr                ), //o
    .io_mem_cmd_payload_uncached            (dataCache_1_io_mem_cmd_payload_uncached          ), //o
    .io_mem_cmd_payload_address             (dataCache_1_io_mem_cmd_payload_address[31:0]     ), //o
    .io_mem_cmd_payload_data                (dataCache_1_io_mem_cmd_payload_data[31:0]        ), //o
    .io_mem_cmd_payload_mask                (dataCache_1_io_mem_cmd_payload_mask[3:0]         ), //o
    .io_mem_cmd_payload_size                (dataCache_1_io_mem_cmd_payload_size[2:0]         ), //o
    .io_mem_cmd_payload_last                (dataCache_1_io_mem_cmd_payload_last              ), //o
    .io_mem_rsp_valid                       (dBus_rsp_valid                                   ), //i
    .io_mem_rsp_payload_last                (dBus_rsp_payload_last                            ), //i
    .io_mem_rsp_payload_data                (dBus_rsp_payload_data[31:0]                      ), //i
    .io_mem_rsp_payload_error               (dBus_rsp_payload_error                           ), //i
    .clk                                    (clk                                              ), //i
    .reset                                  (reset                                            )  //i
  );
  always @(*) begin
    case(_zz_IBusCachedPlugin_jump_pcLoad_payload_6)
      2'b00 : _zz_IBusCachedPlugin_jump_pcLoad_payload_5 = DBusCachedPlugin_redoBranch_payload;
      2'b01 : _zz_IBusCachedPlugin_jump_pcLoad_payload_5 = CsrPlugin_jumpInterface_payload;
      2'b10 : _zz_IBusCachedPlugin_jump_pcLoad_payload_5 = BranchPlugin_jumpInterface_payload;
      default : _zz_IBusCachedPlugin_jump_pcLoad_payload_5 = IBusCachedPlugin_predictionJumpInterface_payload;
    endcase
  end

  always @(*) begin
    case(_zz_writeBack_DBusCachedPlugin_rspShifted_1)
      2'b00 : _zz_writeBack_DBusCachedPlugin_rspShifted = writeBack_DBusCachedPlugin_rspSplits_0;
      2'b01 : _zz_writeBack_DBusCachedPlugin_rspShifted = writeBack_DBusCachedPlugin_rspSplits_1;
      2'b10 : _zz_writeBack_DBusCachedPlugin_rspShifted = writeBack_DBusCachedPlugin_rspSplits_2;
      default : _zz_writeBack_DBusCachedPlugin_rspShifted = writeBack_DBusCachedPlugin_rspSplits_3;
    endcase
  end

  always @(*) begin
    case(_zz_writeBack_DBusCachedPlugin_rspShifted_3)
      1'b0 : _zz_writeBack_DBusCachedPlugin_rspShifted_2 = writeBack_DBusCachedPlugin_rspSplits_1;
      default : _zz_writeBack_DBusCachedPlugin_rspShifted_2 = writeBack_DBusCachedPlugin_rspSplits_3;
    endcase
  end

  always @(*) begin
    case(execute_PmpPlugin_fsm_fsmCounter)
      4'b0000 : _zz_when_PmpPlugin_l246 = PmpPlugin_pmpcfg_0;
      4'b0001 : _zz_when_PmpPlugin_l246 = PmpPlugin_pmpcfg_1;
      4'b0010 : _zz_when_PmpPlugin_l246 = PmpPlugin_pmpcfg_2;
      4'b0011 : _zz_when_PmpPlugin_l246 = PmpPlugin_pmpcfg_3;
      4'b0100 : _zz_when_PmpPlugin_l246 = PmpPlugin_pmpcfg_4;
      4'b0101 : _zz_when_PmpPlugin_l246 = PmpPlugin_pmpcfg_5;
      4'b0110 : _zz_when_PmpPlugin_l246 = PmpPlugin_pmpcfg_6;
      4'b0111 : _zz_when_PmpPlugin_l246 = PmpPlugin_pmpcfg_7;
      4'b1000 : _zz_when_PmpPlugin_l246 = PmpPlugin_pmpcfg_8;
      4'b1001 : _zz_when_PmpPlugin_l246 = PmpPlugin_pmpcfg_9;
      4'b1010 : _zz_when_PmpPlugin_l246 = PmpPlugin_pmpcfg_10;
      4'b1011 : _zz_when_PmpPlugin_l246 = PmpPlugin_pmpcfg_11;
      4'b1100 : _zz_when_PmpPlugin_l246 = PmpPlugin_pmpcfg_12;
      4'b1101 : _zz_when_PmpPlugin_l246 = PmpPlugin_pmpcfg_13;
      4'b1110 : _zz_when_PmpPlugin_l246 = PmpPlugin_pmpcfg_14;
      default : _zz_when_PmpPlugin_l246 = PmpPlugin_pmpcfg_15;
    endcase
  end

  always @(*) begin
    case(_zz_PmpPlugin_dGuard_hits_0_2)
      4'b0000 : _zz_PmpPlugin_dGuard_hits_0_1 = PmpPlugin_mask_0;
      4'b0001 : _zz_PmpPlugin_dGuard_hits_0_1 = PmpPlugin_mask_1;
      4'b0010 : _zz_PmpPlugin_dGuard_hits_0_1 = PmpPlugin_mask_2;
      4'b0011 : _zz_PmpPlugin_dGuard_hits_0_1 = PmpPlugin_mask_3;
      4'b0100 : _zz_PmpPlugin_dGuard_hits_0_1 = PmpPlugin_mask_4;
      4'b0101 : _zz_PmpPlugin_dGuard_hits_0_1 = PmpPlugin_mask_5;
      4'b0110 : _zz_PmpPlugin_dGuard_hits_0_1 = PmpPlugin_mask_6;
      4'b0111 : _zz_PmpPlugin_dGuard_hits_0_1 = PmpPlugin_mask_7;
      4'b1000 : _zz_PmpPlugin_dGuard_hits_0_1 = PmpPlugin_mask_8;
      4'b1001 : _zz_PmpPlugin_dGuard_hits_0_1 = PmpPlugin_mask_9;
      4'b1010 : _zz_PmpPlugin_dGuard_hits_0_1 = PmpPlugin_mask_10;
      4'b1011 : _zz_PmpPlugin_dGuard_hits_0_1 = PmpPlugin_mask_11;
      4'b1100 : _zz_PmpPlugin_dGuard_hits_0_1 = PmpPlugin_mask_12;
      4'b1101 : _zz_PmpPlugin_dGuard_hits_0_1 = PmpPlugin_mask_13;
      4'b1110 : _zz_PmpPlugin_dGuard_hits_0_1 = PmpPlugin_mask_14;
      default : _zz_PmpPlugin_dGuard_hits_0_1 = PmpPlugin_mask_15;
    endcase
  end

  always @(*) begin
    case(_zz_PmpPlugin_dGuard_hits_0_4)
      4'b0000 : _zz_PmpPlugin_dGuard_hits_0_3 = PmpPlugin_base_0;
      4'b0001 : _zz_PmpPlugin_dGuard_hits_0_3 = PmpPlugin_base_1;
      4'b0010 : _zz_PmpPlugin_dGuard_hits_0_3 = PmpPlugin_base_2;
      4'b0011 : _zz_PmpPlugin_dGuard_hits_0_3 = PmpPlugin_base_3;
      4'b0100 : _zz_PmpPlugin_dGuard_hits_0_3 = PmpPlugin_base_4;
      4'b0101 : _zz_PmpPlugin_dGuard_hits_0_3 = PmpPlugin_base_5;
      4'b0110 : _zz_PmpPlugin_dGuard_hits_0_3 = PmpPlugin_base_6;
      4'b0111 : _zz_PmpPlugin_dGuard_hits_0_3 = PmpPlugin_base_7;
      4'b1000 : _zz_PmpPlugin_dGuard_hits_0_3 = PmpPlugin_base_8;
      4'b1001 : _zz_PmpPlugin_dGuard_hits_0_3 = PmpPlugin_base_9;
      4'b1010 : _zz_PmpPlugin_dGuard_hits_0_3 = PmpPlugin_base_10;
      4'b1011 : _zz_PmpPlugin_dGuard_hits_0_3 = PmpPlugin_base_11;
      4'b1100 : _zz_PmpPlugin_dGuard_hits_0_3 = PmpPlugin_base_12;
      4'b1101 : _zz_PmpPlugin_dGuard_hits_0_3 = PmpPlugin_base_13;
      4'b1110 : _zz_PmpPlugin_dGuard_hits_0_3 = PmpPlugin_base_14;
      default : _zz_PmpPlugin_dGuard_hits_0_3 = PmpPlugin_base_15;
    endcase
  end

  always @(*) begin
    case(_zz_PmpPlugin_dGuard_hits_1_1)
      4'b0000 : _zz_PmpPlugin_dGuard_hits_1 = PmpPlugin_mask_0;
      4'b0001 : _zz_PmpPlugin_dGuard_hits_1 = PmpPlugin_mask_1;
      4'b0010 : _zz_PmpPlugin_dGuard_hits_1 = PmpPlugin_mask_2;
      4'b0011 : _zz_PmpPlugin_dGuard_hits_1 = PmpPlugin_mask_3;
      4'b0100 : _zz_PmpPlugin_dGuard_hits_1 = PmpPlugin_mask_4;
      4'b0101 : _zz_PmpPlugin_dGuard_hits_1 = PmpPlugin_mask_5;
      4'b0110 : _zz_PmpPlugin_dGuard_hits_1 = PmpPlugin_mask_6;
      4'b0111 : _zz_PmpPlugin_dGuard_hits_1 = PmpPlugin_mask_7;
      4'b1000 : _zz_PmpPlugin_dGuard_hits_1 = PmpPlugin_mask_8;
      4'b1001 : _zz_PmpPlugin_dGuard_hits_1 = PmpPlugin_mask_9;
      4'b1010 : _zz_PmpPlugin_dGuard_hits_1 = PmpPlugin_mask_10;
      4'b1011 : _zz_PmpPlugin_dGuard_hits_1 = PmpPlugin_mask_11;
      4'b1100 : _zz_PmpPlugin_dGuard_hits_1 = PmpPlugin_mask_12;
      4'b1101 : _zz_PmpPlugin_dGuard_hits_1 = PmpPlugin_mask_13;
      4'b1110 : _zz_PmpPlugin_dGuard_hits_1 = PmpPlugin_mask_14;
      default : _zz_PmpPlugin_dGuard_hits_1 = PmpPlugin_mask_15;
    endcase
  end

  always @(*) begin
    case(_zz_PmpPlugin_dGuard_hits_1_3)
      4'b0000 : _zz_PmpPlugin_dGuard_hits_1_2 = PmpPlugin_base_0;
      4'b0001 : _zz_PmpPlugin_dGuard_hits_1_2 = PmpPlugin_base_1;
      4'b0010 : _zz_PmpPlugin_dGuard_hits_1_2 = PmpPlugin_base_2;
      4'b0011 : _zz_PmpPlugin_dGuard_hits_1_2 = PmpPlugin_base_3;
      4'b0100 : _zz_PmpPlugin_dGuard_hits_1_2 = PmpPlugin_base_4;
      4'b0101 : _zz_PmpPlugin_dGuard_hits_1_2 = PmpPlugin_base_5;
      4'b0110 : _zz_PmpPlugin_dGuard_hits_1_2 = PmpPlugin_base_6;
      4'b0111 : _zz_PmpPlugin_dGuard_hits_1_2 = PmpPlugin_base_7;
      4'b1000 : _zz_PmpPlugin_dGuard_hits_1_2 = PmpPlugin_base_8;
      4'b1001 : _zz_PmpPlugin_dGuard_hits_1_2 = PmpPlugin_base_9;
      4'b1010 : _zz_PmpPlugin_dGuard_hits_1_2 = PmpPlugin_base_10;
      4'b1011 : _zz_PmpPlugin_dGuard_hits_1_2 = PmpPlugin_base_11;
      4'b1100 : _zz_PmpPlugin_dGuard_hits_1_2 = PmpPlugin_base_12;
      4'b1101 : _zz_PmpPlugin_dGuard_hits_1_2 = PmpPlugin_base_13;
      4'b1110 : _zz_PmpPlugin_dGuard_hits_1_2 = PmpPlugin_base_14;
      default : _zz_PmpPlugin_dGuard_hits_1_2 = PmpPlugin_base_15;
    endcase
  end

  always @(*) begin
    case(_zz_PmpPlugin_dGuard_hits_2_1)
      4'b0000 : _zz_PmpPlugin_dGuard_hits_2 = PmpPlugin_mask_0;
      4'b0001 : _zz_PmpPlugin_dGuard_hits_2 = PmpPlugin_mask_1;
      4'b0010 : _zz_PmpPlugin_dGuard_hits_2 = PmpPlugin_mask_2;
      4'b0011 : _zz_PmpPlugin_dGuard_hits_2 = PmpPlugin_mask_3;
      4'b0100 : _zz_PmpPlugin_dGuard_hits_2 = PmpPlugin_mask_4;
      4'b0101 : _zz_PmpPlugin_dGuard_hits_2 = PmpPlugin_mask_5;
      4'b0110 : _zz_PmpPlugin_dGuard_hits_2 = PmpPlugin_mask_6;
      4'b0111 : _zz_PmpPlugin_dGuard_hits_2 = PmpPlugin_mask_7;
      4'b1000 : _zz_PmpPlugin_dGuard_hits_2 = PmpPlugin_mask_8;
      4'b1001 : _zz_PmpPlugin_dGuard_hits_2 = PmpPlugin_mask_9;
      4'b1010 : _zz_PmpPlugin_dGuard_hits_2 = PmpPlugin_mask_10;
      4'b1011 : _zz_PmpPlugin_dGuard_hits_2 = PmpPlugin_mask_11;
      4'b1100 : _zz_PmpPlugin_dGuard_hits_2 = PmpPlugin_mask_12;
      4'b1101 : _zz_PmpPlugin_dGuard_hits_2 = PmpPlugin_mask_13;
      4'b1110 : _zz_PmpPlugin_dGuard_hits_2 = PmpPlugin_mask_14;
      default : _zz_PmpPlugin_dGuard_hits_2 = PmpPlugin_mask_15;
    endcase
  end

  always @(*) begin
    case(_zz_PmpPlugin_dGuard_hits_2_3)
      4'b0000 : _zz_PmpPlugin_dGuard_hits_2_2 = PmpPlugin_base_0;
      4'b0001 : _zz_PmpPlugin_dGuard_hits_2_2 = PmpPlugin_base_1;
      4'b0010 : _zz_PmpPlugin_dGuard_hits_2_2 = PmpPlugin_base_2;
      4'b0011 : _zz_PmpPlugin_dGuard_hits_2_2 = PmpPlugin_base_3;
      4'b0100 : _zz_PmpPlugin_dGuard_hits_2_2 = PmpPlugin_base_4;
      4'b0101 : _zz_PmpPlugin_dGuard_hits_2_2 = PmpPlugin_base_5;
      4'b0110 : _zz_PmpPlugin_dGuard_hits_2_2 = PmpPlugin_base_6;
      4'b0111 : _zz_PmpPlugin_dGuard_hits_2_2 = PmpPlugin_base_7;
      4'b1000 : _zz_PmpPlugin_dGuard_hits_2_2 = PmpPlugin_base_8;
      4'b1001 : _zz_PmpPlugin_dGuard_hits_2_2 = PmpPlugin_base_9;
      4'b1010 : _zz_PmpPlugin_dGuard_hits_2_2 = PmpPlugin_base_10;
      4'b1011 : _zz_PmpPlugin_dGuard_hits_2_2 = PmpPlugin_base_11;
      4'b1100 : _zz_PmpPlugin_dGuard_hits_2_2 = PmpPlugin_base_12;
      4'b1101 : _zz_PmpPlugin_dGuard_hits_2_2 = PmpPlugin_base_13;
      4'b1110 : _zz_PmpPlugin_dGuard_hits_2_2 = PmpPlugin_base_14;
      default : _zz_PmpPlugin_dGuard_hits_2_2 = PmpPlugin_base_15;
    endcase
  end

  always @(*) begin
    case(_zz_PmpPlugin_dGuard_hits_3_1)
      4'b0000 : _zz_PmpPlugin_dGuard_hits_3 = PmpPlugin_mask_0;
      4'b0001 : _zz_PmpPlugin_dGuard_hits_3 = PmpPlugin_mask_1;
      4'b0010 : _zz_PmpPlugin_dGuard_hits_3 = PmpPlugin_mask_2;
      4'b0011 : _zz_PmpPlugin_dGuard_hits_3 = PmpPlugin_mask_3;
      4'b0100 : _zz_PmpPlugin_dGuard_hits_3 = PmpPlugin_mask_4;
      4'b0101 : _zz_PmpPlugin_dGuard_hits_3 = PmpPlugin_mask_5;
      4'b0110 : _zz_PmpPlugin_dGuard_hits_3 = PmpPlugin_mask_6;
      4'b0111 : _zz_PmpPlugin_dGuard_hits_3 = PmpPlugin_mask_7;
      4'b1000 : _zz_PmpPlugin_dGuard_hits_3 = PmpPlugin_mask_8;
      4'b1001 : _zz_PmpPlugin_dGuard_hits_3 = PmpPlugin_mask_9;
      4'b1010 : _zz_PmpPlugin_dGuard_hits_3 = PmpPlugin_mask_10;
      4'b1011 : _zz_PmpPlugin_dGuard_hits_3 = PmpPlugin_mask_11;
      4'b1100 : _zz_PmpPlugin_dGuard_hits_3 = PmpPlugin_mask_12;
      4'b1101 : _zz_PmpPlugin_dGuard_hits_3 = PmpPlugin_mask_13;
      4'b1110 : _zz_PmpPlugin_dGuard_hits_3 = PmpPlugin_mask_14;
      default : _zz_PmpPlugin_dGuard_hits_3 = PmpPlugin_mask_15;
    endcase
  end

  always @(*) begin
    case(_zz_PmpPlugin_dGuard_hits_3_3)
      4'b0000 : _zz_PmpPlugin_dGuard_hits_3_2 = PmpPlugin_base_0;
      4'b0001 : _zz_PmpPlugin_dGuard_hits_3_2 = PmpPlugin_base_1;
      4'b0010 : _zz_PmpPlugin_dGuard_hits_3_2 = PmpPlugin_base_2;
      4'b0011 : _zz_PmpPlugin_dGuard_hits_3_2 = PmpPlugin_base_3;
      4'b0100 : _zz_PmpPlugin_dGuard_hits_3_2 = PmpPlugin_base_4;
      4'b0101 : _zz_PmpPlugin_dGuard_hits_3_2 = PmpPlugin_base_5;
      4'b0110 : _zz_PmpPlugin_dGuard_hits_3_2 = PmpPlugin_base_6;
      4'b0111 : _zz_PmpPlugin_dGuard_hits_3_2 = PmpPlugin_base_7;
      4'b1000 : _zz_PmpPlugin_dGuard_hits_3_2 = PmpPlugin_base_8;
      4'b1001 : _zz_PmpPlugin_dGuard_hits_3_2 = PmpPlugin_base_9;
      4'b1010 : _zz_PmpPlugin_dGuard_hits_3_2 = PmpPlugin_base_10;
      4'b1011 : _zz_PmpPlugin_dGuard_hits_3_2 = PmpPlugin_base_11;
      4'b1100 : _zz_PmpPlugin_dGuard_hits_3_2 = PmpPlugin_base_12;
      4'b1101 : _zz_PmpPlugin_dGuard_hits_3_2 = PmpPlugin_base_13;
      4'b1110 : _zz_PmpPlugin_dGuard_hits_3_2 = PmpPlugin_base_14;
      default : _zz_PmpPlugin_dGuard_hits_3_2 = PmpPlugin_base_15;
    endcase
  end

  always @(*) begin
    case(_zz_PmpPlugin_dGuard_hits_4_1)
      4'b0000 : _zz_PmpPlugin_dGuard_hits_4 = PmpPlugin_mask_0;
      4'b0001 : _zz_PmpPlugin_dGuard_hits_4 = PmpPlugin_mask_1;
      4'b0010 : _zz_PmpPlugin_dGuard_hits_4 = PmpPlugin_mask_2;
      4'b0011 : _zz_PmpPlugin_dGuard_hits_4 = PmpPlugin_mask_3;
      4'b0100 : _zz_PmpPlugin_dGuard_hits_4 = PmpPlugin_mask_4;
      4'b0101 : _zz_PmpPlugin_dGuard_hits_4 = PmpPlugin_mask_5;
      4'b0110 : _zz_PmpPlugin_dGuard_hits_4 = PmpPlugin_mask_6;
      4'b0111 : _zz_PmpPlugin_dGuard_hits_4 = PmpPlugin_mask_7;
      4'b1000 : _zz_PmpPlugin_dGuard_hits_4 = PmpPlugin_mask_8;
      4'b1001 : _zz_PmpPlugin_dGuard_hits_4 = PmpPlugin_mask_9;
      4'b1010 : _zz_PmpPlugin_dGuard_hits_4 = PmpPlugin_mask_10;
      4'b1011 : _zz_PmpPlugin_dGuard_hits_4 = PmpPlugin_mask_11;
      4'b1100 : _zz_PmpPlugin_dGuard_hits_4 = PmpPlugin_mask_12;
      4'b1101 : _zz_PmpPlugin_dGuard_hits_4 = PmpPlugin_mask_13;
      4'b1110 : _zz_PmpPlugin_dGuard_hits_4 = PmpPlugin_mask_14;
      default : _zz_PmpPlugin_dGuard_hits_4 = PmpPlugin_mask_15;
    endcase
  end

  always @(*) begin
    case(_zz_PmpPlugin_dGuard_hits_4_3)
      4'b0000 : _zz_PmpPlugin_dGuard_hits_4_2 = PmpPlugin_base_0;
      4'b0001 : _zz_PmpPlugin_dGuard_hits_4_2 = PmpPlugin_base_1;
      4'b0010 : _zz_PmpPlugin_dGuard_hits_4_2 = PmpPlugin_base_2;
      4'b0011 : _zz_PmpPlugin_dGuard_hits_4_2 = PmpPlugin_base_3;
      4'b0100 : _zz_PmpPlugin_dGuard_hits_4_2 = PmpPlugin_base_4;
      4'b0101 : _zz_PmpPlugin_dGuard_hits_4_2 = PmpPlugin_base_5;
      4'b0110 : _zz_PmpPlugin_dGuard_hits_4_2 = PmpPlugin_base_6;
      4'b0111 : _zz_PmpPlugin_dGuard_hits_4_2 = PmpPlugin_base_7;
      4'b1000 : _zz_PmpPlugin_dGuard_hits_4_2 = PmpPlugin_base_8;
      4'b1001 : _zz_PmpPlugin_dGuard_hits_4_2 = PmpPlugin_base_9;
      4'b1010 : _zz_PmpPlugin_dGuard_hits_4_2 = PmpPlugin_base_10;
      4'b1011 : _zz_PmpPlugin_dGuard_hits_4_2 = PmpPlugin_base_11;
      4'b1100 : _zz_PmpPlugin_dGuard_hits_4_2 = PmpPlugin_base_12;
      4'b1101 : _zz_PmpPlugin_dGuard_hits_4_2 = PmpPlugin_base_13;
      4'b1110 : _zz_PmpPlugin_dGuard_hits_4_2 = PmpPlugin_base_14;
      default : _zz_PmpPlugin_dGuard_hits_4_2 = PmpPlugin_base_15;
    endcase
  end

  always @(*) begin
    case(_zz_PmpPlugin_dGuard_hits_5_1)
      4'b0000 : _zz_PmpPlugin_dGuard_hits_5 = PmpPlugin_mask_0;
      4'b0001 : _zz_PmpPlugin_dGuard_hits_5 = PmpPlugin_mask_1;
      4'b0010 : _zz_PmpPlugin_dGuard_hits_5 = PmpPlugin_mask_2;
      4'b0011 : _zz_PmpPlugin_dGuard_hits_5 = PmpPlugin_mask_3;
      4'b0100 : _zz_PmpPlugin_dGuard_hits_5 = PmpPlugin_mask_4;
      4'b0101 : _zz_PmpPlugin_dGuard_hits_5 = PmpPlugin_mask_5;
      4'b0110 : _zz_PmpPlugin_dGuard_hits_5 = PmpPlugin_mask_6;
      4'b0111 : _zz_PmpPlugin_dGuard_hits_5 = PmpPlugin_mask_7;
      4'b1000 : _zz_PmpPlugin_dGuard_hits_5 = PmpPlugin_mask_8;
      4'b1001 : _zz_PmpPlugin_dGuard_hits_5 = PmpPlugin_mask_9;
      4'b1010 : _zz_PmpPlugin_dGuard_hits_5 = PmpPlugin_mask_10;
      4'b1011 : _zz_PmpPlugin_dGuard_hits_5 = PmpPlugin_mask_11;
      4'b1100 : _zz_PmpPlugin_dGuard_hits_5 = PmpPlugin_mask_12;
      4'b1101 : _zz_PmpPlugin_dGuard_hits_5 = PmpPlugin_mask_13;
      4'b1110 : _zz_PmpPlugin_dGuard_hits_5 = PmpPlugin_mask_14;
      default : _zz_PmpPlugin_dGuard_hits_5 = PmpPlugin_mask_15;
    endcase
  end

  always @(*) begin
    case(_zz_PmpPlugin_dGuard_hits_5_3)
      4'b0000 : _zz_PmpPlugin_dGuard_hits_5_2 = PmpPlugin_base_0;
      4'b0001 : _zz_PmpPlugin_dGuard_hits_5_2 = PmpPlugin_base_1;
      4'b0010 : _zz_PmpPlugin_dGuard_hits_5_2 = PmpPlugin_base_2;
      4'b0011 : _zz_PmpPlugin_dGuard_hits_5_2 = PmpPlugin_base_3;
      4'b0100 : _zz_PmpPlugin_dGuard_hits_5_2 = PmpPlugin_base_4;
      4'b0101 : _zz_PmpPlugin_dGuard_hits_5_2 = PmpPlugin_base_5;
      4'b0110 : _zz_PmpPlugin_dGuard_hits_5_2 = PmpPlugin_base_6;
      4'b0111 : _zz_PmpPlugin_dGuard_hits_5_2 = PmpPlugin_base_7;
      4'b1000 : _zz_PmpPlugin_dGuard_hits_5_2 = PmpPlugin_base_8;
      4'b1001 : _zz_PmpPlugin_dGuard_hits_5_2 = PmpPlugin_base_9;
      4'b1010 : _zz_PmpPlugin_dGuard_hits_5_2 = PmpPlugin_base_10;
      4'b1011 : _zz_PmpPlugin_dGuard_hits_5_2 = PmpPlugin_base_11;
      4'b1100 : _zz_PmpPlugin_dGuard_hits_5_2 = PmpPlugin_base_12;
      4'b1101 : _zz_PmpPlugin_dGuard_hits_5_2 = PmpPlugin_base_13;
      4'b1110 : _zz_PmpPlugin_dGuard_hits_5_2 = PmpPlugin_base_14;
      default : _zz_PmpPlugin_dGuard_hits_5_2 = PmpPlugin_base_15;
    endcase
  end

  always @(*) begin
    case(_zz_PmpPlugin_dGuard_hits_6_1)
      4'b0000 : _zz_PmpPlugin_dGuard_hits_6 = PmpPlugin_mask_0;
      4'b0001 : _zz_PmpPlugin_dGuard_hits_6 = PmpPlugin_mask_1;
      4'b0010 : _zz_PmpPlugin_dGuard_hits_6 = PmpPlugin_mask_2;
      4'b0011 : _zz_PmpPlugin_dGuard_hits_6 = PmpPlugin_mask_3;
      4'b0100 : _zz_PmpPlugin_dGuard_hits_6 = PmpPlugin_mask_4;
      4'b0101 : _zz_PmpPlugin_dGuard_hits_6 = PmpPlugin_mask_5;
      4'b0110 : _zz_PmpPlugin_dGuard_hits_6 = PmpPlugin_mask_6;
      4'b0111 : _zz_PmpPlugin_dGuard_hits_6 = PmpPlugin_mask_7;
      4'b1000 : _zz_PmpPlugin_dGuard_hits_6 = PmpPlugin_mask_8;
      4'b1001 : _zz_PmpPlugin_dGuard_hits_6 = PmpPlugin_mask_9;
      4'b1010 : _zz_PmpPlugin_dGuard_hits_6 = PmpPlugin_mask_10;
      4'b1011 : _zz_PmpPlugin_dGuard_hits_6 = PmpPlugin_mask_11;
      4'b1100 : _zz_PmpPlugin_dGuard_hits_6 = PmpPlugin_mask_12;
      4'b1101 : _zz_PmpPlugin_dGuard_hits_6 = PmpPlugin_mask_13;
      4'b1110 : _zz_PmpPlugin_dGuard_hits_6 = PmpPlugin_mask_14;
      default : _zz_PmpPlugin_dGuard_hits_6 = PmpPlugin_mask_15;
    endcase
  end

  always @(*) begin
    case(_zz_PmpPlugin_dGuard_hits_6_3)
      4'b0000 : _zz_PmpPlugin_dGuard_hits_6_2 = PmpPlugin_base_0;
      4'b0001 : _zz_PmpPlugin_dGuard_hits_6_2 = PmpPlugin_base_1;
      4'b0010 : _zz_PmpPlugin_dGuard_hits_6_2 = PmpPlugin_base_2;
      4'b0011 : _zz_PmpPlugin_dGuard_hits_6_2 = PmpPlugin_base_3;
      4'b0100 : _zz_PmpPlugin_dGuard_hits_6_2 = PmpPlugin_base_4;
      4'b0101 : _zz_PmpPlugin_dGuard_hits_6_2 = PmpPlugin_base_5;
      4'b0110 : _zz_PmpPlugin_dGuard_hits_6_2 = PmpPlugin_base_6;
      4'b0111 : _zz_PmpPlugin_dGuard_hits_6_2 = PmpPlugin_base_7;
      4'b1000 : _zz_PmpPlugin_dGuard_hits_6_2 = PmpPlugin_base_8;
      4'b1001 : _zz_PmpPlugin_dGuard_hits_6_2 = PmpPlugin_base_9;
      4'b1010 : _zz_PmpPlugin_dGuard_hits_6_2 = PmpPlugin_base_10;
      4'b1011 : _zz_PmpPlugin_dGuard_hits_6_2 = PmpPlugin_base_11;
      4'b1100 : _zz_PmpPlugin_dGuard_hits_6_2 = PmpPlugin_base_12;
      4'b1101 : _zz_PmpPlugin_dGuard_hits_6_2 = PmpPlugin_base_13;
      4'b1110 : _zz_PmpPlugin_dGuard_hits_6_2 = PmpPlugin_base_14;
      default : _zz_PmpPlugin_dGuard_hits_6_2 = PmpPlugin_base_15;
    endcase
  end

  always @(*) begin
    case(_zz_PmpPlugin_dGuard_hits_7_1)
      4'b0000 : _zz_PmpPlugin_dGuard_hits_7 = PmpPlugin_mask_0;
      4'b0001 : _zz_PmpPlugin_dGuard_hits_7 = PmpPlugin_mask_1;
      4'b0010 : _zz_PmpPlugin_dGuard_hits_7 = PmpPlugin_mask_2;
      4'b0011 : _zz_PmpPlugin_dGuard_hits_7 = PmpPlugin_mask_3;
      4'b0100 : _zz_PmpPlugin_dGuard_hits_7 = PmpPlugin_mask_4;
      4'b0101 : _zz_PmpPlugin_dGuard_hits_7 = PmpPlugin_mask_5;
      4'b0110 : _zz_PmpPlugin_dGuard_hits_7 = PmpPlugin_mask_6;
      4'b0111 : _zz_PmpPlugin_dGuard_hits_7 = PmpPlugin_mask_7;
      4'b1000 : _zz_PmpPlugin_dGuard_hits_7 = PmpPlugin_mask_8;
      4'b1001 : _zz_PmpPlugin_dGuard_hits_7 = PmpPlugin_mask_9;
      4'b1010 : _zz_PmpPlugin_dGuard_hits_7 = PmpPlugin_mask_10;
      4'b1011 : _zz_PmpPlugin_dGuard_hits_7 = PmpPlugin_mask_11;
      4'b1100 : _zz_PmpPlugin_dGuard_hits_7 = PmpPlugin_mask_12;
      4'b1101 : _zz_PmpPlugin_dGuard_hits_7 = PmpPlugin_mask_13;
      4'b1110 : _zz_PmpPlugin_dGuard_hits_7 = PmpPlugin_mask_14;
      default : _zz_PmpPlugin_dGuard_hits_7 = PmpPlugin_mask_15;
    endcase
  end

  always @(*) begin
    case(_zz_PmpPlugin_dGuard_hits_7_3)
      4'b0000 : _zz_PmpPlugin_dGuard_hits_7_2 = PmpPlugin_base_0;
      4'b0001 : _zz_PmpPlugin_dGuard_hits_7_2 = PmpPlugin_base_1;
      4'b0010 : _zz_PmpPlugin_dGuard_hits_7_2 = PmpPlugin_base_2;
      4'b0011 : _zz_PmpPlugin_dGuard_hits_7_2 = PmpPlugin_base_3;
      4'b0100 : _zz_PmpPlugin_dGuard_hits_7_2 = PmpPlugin_base_4;
      4'b0101 : _zz_PmpPlugin_dGuard_hits_7_2 = PmpPlugin_base_5;
      4'b0110 : _zz_PmpPlugin_dGuard_hits_7_2 = PmpPlugin_base_6;
      4'b0111 : _zz_PmpPlugin_dGuard_hits_7_2 = PmpPlugin_base_7;
      4'b1000 : _zz_PmpPlugin_dGuard_hits_7_2 = PmpPlugin_base_8;
      4'b1001 : _zz_PmpPlugin_dGuard_hits_7_2 = PmpPlugin_base_9;
      4'b1010 : _zz_PmpPlugin_dGuard_hits_7_2 = PmpPlugin_base_10;
      4'b1011 : _zz_PmpPlugin_dGuard_hits_7_2 = PmpPlugin_base_11;
      4'b1100 : _zz_PmpPlugin_dGuard_hits_7_2 = PmpPlugin_base_12;
      4'b1101 : _zz_PmpPlugin_dGuard_hits_7_2 = PmpPlugin_base_13;
      4'b1110 : _zz_PmpPlugin_dGuard_hits_7_2 = PmpPlugin_base_14;
      default : _zz_PmpPlugin_dGuard_hits_7_2 = PmpPlugin_base_15;
    endcase
  end

  always @(*) begin
    case(_zz_PmpPlugin_dGuard_hits_8_1)
      4'b0000 : _zz_PmpPlugin_dGuard_hits_8 = PmpPlugin_mask_0;
      4'b0001 : _zz_PmpPlugin_dGuard_hits_8 = PmpPlugin_mask_1;
      4'b0010 : _zz_PmpPlugin_dGuard_hits_8 = PmpPlugin_mask_2;
      4'b0011 : _zz_PmpPlugin_dGuard_hits_8 = PmpPlugin_mask_3;
      4'b0100 : _zz_PmpPlugin_dGuard_hits_8 = PmpPlugin_mask_4;
      4'b0101 : _zz_PmpPlugin_dGuard_hits_8 = PmpPlugin_mask_5;
      4'b0110 : _zz_PmpPlugin_dGuard_hits_8 = PmpPlugin_mask_6;
      4'b0111 : _zz_PmpPlugin_dGuard_hits_8 = PmpPlugin_mask_7;
      4'b1000 : _zz_PmpPlugin_dGuard_hits_8 = PmpPlugin_mask_8;
      4'b1001 : _zz_PmpPlugin_dGuard_hits_8 = PmpPlugin_mask_9;
      4'b1010 : _zz_PmpPlugin_dGuard_hits_8 = PmpPlugin_mask_10;
      4'b1011 : _zz_PmpPlugin_dGuard_hits_8 = PmpPlugin_mask_11;
      4'b1100 : _zz_PmpPlugin_dGuard_hits_8 = PmpPlugin_mask_12;
      4'b1101 : _zz_PmpPlugin_dGuard_hits_8 = PmpPlugin_mask_13;
      4'b1110 : _zz_PmpPlugin_dGuard_hits_8 = PmpPlugin_mask_14;
      default : _zz_PmpPlugin_dGuard_hits_8 = PmpPlugin_mask_15;
    endcase
  end

  always @(*) begin
    case(_zz_PmpPlugin_dGuard_hits_8_3)
      4'b0000 : _zz_PmpPlugin_dGuard_hits_8_2 = PmpPlugin_base_0;
      4'b0001 : _zz_PmpPlugin_dGuard_hits_8_2 = PmpPlugin_base_1;
      4'b0010 : _zz_PmpPlugin_dGuard_hits_8_2 = PmpPlugin_base_2;
      4'b0011 : _zz_PmpPlugin_dGuard_hits_8_2 = PmpPlugin_base_3;
      4'b0100 : _zz_PmpPlugin_dGuard_hits_8_2 = PmpPlugin_base_4;
      4'b0101 : _zz_PmpPlugin_dGuard_hits_8_2 = PmpPlugin_base_5;
      4'b0110 : _zz_PmpPlugin_dGuard_hits_8_2 = PmpPlugin_base_6;
      4'b0111 : _zz_PmpPlugin_dGuard_hits_8_2 = PmpPlugin_base_7;
      4'b1000 : _zz_PmpPlugin_dGuard_hits_8_2 = PmpPlugin_base_8;
      4'b1001 : _zz_PmpPlugin_dGuard_hits_8_2 = PmpPlugin_base_9;
      4'b1010 : _zz_PmpPlugin_dGuard_hits_8_2 = PmpPlugin_base_10;
      4'b1011 : _zz_PmpPlugin_dGuard_hits_8_2 = PmpPlugin_base_11;
      4'b1100 : _zz_PmpPlugin_dGuard_hits_8_2 = PmpPlugin_base_12;
      4'b1101 : _zz_PmpPlugin_dGuard_hits_8_2 = PmpPlugin_base_13;
      4'b1110 : _zz_PmpPlugin_dGuard_hits_8_2 = PmpPlugin_base_14;
      default : _zz_PmpPlugin_dGuard_hits_8_2 = PmpPlugin_base_15;
    endcase
  end

  always @(*) begin
    case(_zz_PmpPlugin_dGuard_hits_9_1)
      4'b0000 : _zz_PmpPlugin_dGuard_hits_9 = PmpPlugin_mask_0;
      4'b0001 : _zz_PmpPlugin_dGuard_hits_9 = PmpPlugin_mask_1;
      4'b0010 : _zz_PmpPlugin_dGuard_hits_9 = PmpPlugin_mask_2;
      4'b0011 : _zz_PmpPlugin_dGuard_hits_9 = PmpPlugin_mask_3;
      4'b0100 : _zz_PmpPlugin_dGuard_hits_9 = PmpPlugin_mask_4;
      4'b0101 : _zz_PmpPlugin_dGuard_hits_9 = PmpPlugin_mask_5;
      4'b0110 : _zz_PmpPlugin_dGuard_hits_9 = PmpPlugin_mask_6;
      4'b0111 : _zz_PmpPlugin_dGuard_hits_9 = PmpPlugin_mask_7;
      4'b1000 : _zz_PmpPlugin_dGuard_hits_9 = PmpPlugin_mask_8;
      4'b1001 : _zz_PmpPlugin_dGuard_hits_9 = PmpPlugin_mask_9;
      4'b1010 : _zz_PmpPlugin_dGuard_hits_9 = PmpPlugin_mask_10;
      4'b1011 : _zz_PmpPlugin_dGuard_hits_9 = PmpPlugin_mask_11;
      4'b1100 : _zz_PmpPlugin_dGuard_hits_9 = PmpPlugin_mask_12;
      4'b1101 : _zz_PmpPlugin_dGuard_hits_9 = PmpPlugin_mask_13;
      4'b1110 : _zz_PmpPlugin_dGuard_hits_9 = PmpPlugin_mask_14;
      default : _zz_PmpPlugin_dGuard_hits_9 = PmpPlugin_mask_15;
    endcase
  end

  always @(*) begin
    case(_zz_PmpPlugin_dGuard_hits_9_3)
      4'b0000 : _zz_PmpPlugin_dGuard_hits_9_2 = PmpPlugin_base_0;
      4'b0001 : _zz_PmpPlugin_dGuard_hits_9_2 = PmpPlugin_base_1;
      4'b0010 : _zz_PmpPlugin_dGuard_hits_9_2 = PmpPlugin_base_2;
      4'b0011 : _zz_PmpPlugin_dGuard_hits_9_2 = PmpPlugin_base_3;
      4'b0100 : _zz_PmpPlugin_dGuard_hits_9_2 = PmpPlugin_base_4;
      4'b0101 : _zz_PmpPlugin_dGuard_hits_9_2 = PmpPlugin_base_5;
      4'b0110 : _zz_PmpPlugin_dGuard_hits_9_2 = PmpPlugin_base_6;
      4'b0111 : _zz_PmpPlugin_dGuard_hits_9_2 = PmpPlugin_base_7;
      4'b1000 : _zz_PmpPlugin_dGuard_hits_9_2 = PmpPlugin_base_8;
      4'b1001 : _zz_PmpPlugin_dGuard_hits_9_2 = PmpPlugin_base_9;
      4'b1010 : _zz_PmpPlugin_dGuard_hits_9_2 = PmpPlugin_base_10;
      4'b1011 : _zz_PmpPlugin_dGuard_hits_9_2 = PmpPlugin_base_11;
      4'b1100 : _zz_PmpPlugin_dGuard_hits_9_2 = PmpPlugin_base_12;
      4'b1101 : _zz_PmpPlugin_dGuard_hits_9_2 = PmpPlugin_base_13;
      4'b1110 : _zz_PmpPlugin_dGuard_hits_9_2 = PmpPlugin_base_14;
      default : _zz_PmpPlugin_dGuard_hits_9_2 = PmpPlugin_base_15;
    endcase
  end

  always @(*) begin
    case(_zz_PmpPlugin_dGuard_hits_10_1)
      4'b0000 : _zz_PmpPlugin_dGuard_hits_10 = PmpPlugin_mask_0;
      4'b0001 : _zz_PmpPlugin_dGuard_hits_10 = PmpPlugin_mask_1;
      4'b0010 : _zz_PmpPlugin_dGuard_hits_10 = PmpPlugin_mask_2;
      4'b0011 : _zz_PmpPlugin_dGuard_hits_10 = PmpPlugin_mask_3;
      4'b0100 : _zz_PmpPlugin_dGuard_hits_10 = PmpPlugin_mask_4;
      4'b0101 : _zz_PmpPlugin_dGuard_hits_10 = PmpPlugin_mask_5;
      4'b0110 : _zz_PmpPlugin_dGuard_hits_10 = PmpPlugin_mask_6;
      4'b0111 : _zz_PmpPlugin_dGuard_hits_10 = PmpPlugin_mask_7;
      4'b1000 : _zz_PmpPlugin_dGuard_hits_10 = PmpPlugin_mask_8;
      4'b1001 : _zz_PmpPlugin_dGuard_hits_10 = PmpPlugin_mask_9;
      4'b1010 : _zz_PmpPlugin_dGuard_hits_10 = PmpPlugin_mask_10;
      4'b1011 : _zz_PmpPlugin_dGuard_hits_10 = PmpPlugin_mask_11;
      4'b1100 : _zz_PmpPlugin_dGuard_hits_10 = PmpPlugin_mask_12;
      4'b1101 : _zz_PmpPlugin_dGuard_hits_10 = PmpPlugin_mask_13;
      4'b1110 : _zz_PmpPlugin_dGuard_hits_10 = PmpPlugin_mask_14;
      default : _zz_PmpPlugin_dGuard_hits_10 = PmpPlugin_mask_15;
    endcase
  end

  always @(*) begin
    case(_zz_PmpPlugin_dGuard_hits_10_3)
      4'b0000 : _zz_PmpPlugin_dGuard_hits_10_2 = PmpPlugin_base_0;
      4'b0001 : _zz_PmpPlugin_dGuard_hits_10_2 = PmpPlugin_base_1;
      4'b0010 : _zz_PmpPlugin_dGuard_hits_10_2 = PmpPlugin_base_2;
      4'b0011 : _zz_PmpPlugin_dGuard_hits_10_2 = PmpPlugin_base_3;
      4'b0100 : _zz_PmpPlugin_dGuard_hits_10_2 = PmpPlugin_base_4;
      4'b0101 : _zz_PmpPlugin_dGuard_hits_10_2 = PmpPlugin_base_5;
      4'b0110 : _zz_PmpPlugin_dGuard_hits_10_2 = PmpPlugin_base_6;
      4'b0111 : _zz_PmpPlugin_dGuard_hits_10_2 = PmpPlugin_base_7;
      4'b1000 : _zz_PmpPlugin_dGuard_hits_10_2 = PmpPlugin_base_8;
      4'b1001 : _zz_PmpPlugin_dGuard_hits_10_2 = PmpPlugin_base_9;
      4'b1010 : _zz_PmpPlugin_dGuard_hits_10_2 = PmpPlugin_base_10;
      4'b1011 : _zz_PmpPlugin_dGuard_hits_10_2 = PmpPlugin_base_11;
      4'b1100 : _zz_PmpPlugin_dGuard_hits_10_2 = PmpPlugin_base_12;
      4'b1101 : _zz_PmpPlugin_dGuard_hits_10_2 = PmpPlugin_base_13;
      4'b1110 : _zz_PmpPlugin_dGuard_hits_10_2 = PmpPlugin_base_14;
      default : _zz_PmpPlugin_dGuard_hits_10_2 = PmpPlugin_base_15;
    endcase
  end

  always @(*) begin
    case(_zz_PmpPlugin_dGuard_hits_11_1)
      4'b0000 : _zz_PmpPlugin_dGuard_hits_11 = PmpPlugin_mask_0;
      4'b0001 : _zz_PmpPlugin_dGuard_hits_11 = PmpPlugin_mask_1;
      4'b0010 : _zz_PmpPlugin_dGuard_hits_11 = PmpPlugin_mask_2;
      4'b0011 : _zz_PmpPlugin_dGuard_hits_11 = PmpPlugin_mask_3;
      4'b0100 : _zz_PmpPlugin_dGuard_hits_11 = PmpPlugin_mask_4;
      4'b0101 : _zz_PmpPlugin_dGuard_hits_11 = PmpPlugin_mask_5;
      4'b0110 : _zz_PmpPlugin_dGuard_hits_11 = PmpPlugin_mask_6;
      4'b0111 : _zz_PmpPlugin_dGuard_hits_11 = PmpPlugin_mask_7;
      4'b1000 : _zz_PmpPlugin_dGuard_hits_11 = PmpPlugin_mask_8;
      4'b1001 : _zz_PmpPlugin_dGuard_hits_11 = PmpPlugin_mask_9;
      4'b1010 : _zz_PmpPlugin_dGuard_hits_11 = PmpPlugin_mask_10;
      4'b1011 : _zz_PmpPlugin_dGuard_hits_11 = PmpPlugin_mask_11;
      4'b1100 : _zz_PmpPlugin_dGuard_hits_11 = PmpPlugin_mask_12;
      4'b1101 : _zz_PmpPlugin_dGuard_hits_11 = PmpPlugin_mask_13;
      4'b1110 : _zz_PmpPlugin_dGuard_hits_11 = PmpPlugin_mask_14;
      default : _zz_PmpPlugin_dGuard_hits_11 = PmpPlugin_mask_15;
    endcase
  end

  always @(*) begin
    case(_zz_PmpPlugin_dGuard_hits_11_3)
      4'b0000 : _zz_PmpPlugin_dGuard_hits_11_2 = PmpPlugin_base_0;
      4'b0001 : _zz_PmpPlugin_dGuard_hits_11_2 = PmpPlugin_base_1;
      4'b0010 : _zz_PmpPlugin_dGuard_hits_11_2 = PmpPlugin_base_2;
      4'b0011 : _zz_PmpPlugin_dGuard_hits_11_2 = PmpPlugin_base_3;
      4'b0100 : _zz_PmpPlugin_dGuard_hits_11_2 = PmpPlugin_base_4;
      4'b0101 : _zz_PmpPlugin_dGuard_hits_11_2 = PmpPlugin_base_5;
      4'b0110 : _zz_PmpPlugin_dGuard_hits_11_2 = PmpPlugin_base_6;
      4'b0111 : _zz_PmpPlugin_dGuard_hits_11_2 = PmpPlugin_base_7;
      4'b1000 : _zz_PmpPlugin_dGuard_hits_11_2 = PmpPlugin_base_8;
      4'b1001 : _zz_PmpPlugin_dGuard_hits_11_2 = PmpPlugin_base_9;
      4'b1010 : _zz_PmpPlugin_dGuard_hits_11_2 = PmpPlugin_base_10;
      4'b1011 : _zz_PmpPlugin_dGuard_hits_11_2 = PmpPlugin_base_11;
      4'b1100 : _zz_PmpPlugin_dGuard_hits_11_2 = PmpPlugin_base_12;
      4'b1101 : _zz_PmpPlugin_dGuard_hits_11_2 = PmpPlugin_base_13;
      4'b1110 : _zz_PmpPlugin_dGuard_hits_11_2 = PmpPlugin_base_14;
      default : _zz_PmpPlugin_dGuard_hits_11_2 = PmpPlugin_base_15;
    endcase
  end

  always @(*) begin
    case(_zz_PmpPlugin_dGuard_hits_12_1)
      4'b0000 : _zz_PmpPlugin_dGuard_hits_12 = PmpPlugin_mask_0;
      4'b0001 : _zz_PmpPlugin_dGuard_hits_12 = PmpPlugin_mask_1;
      4'b0010 : _zz_PmpPlugin_dGuard_hits_12 = PmpPlugin_mask_2;
      4'b0011 : _zz_PmpPlugin_dGuard_hits_12 = PmpPlugin_mask_3;
      4'b0100 : _zz_PmpPlugin_dGuard_hits_12 = PmpPlugin_mask_4;
      4'b0101 : _zz_PmpPlugin_dGuard_hits_12 = PmpPlugin_mask_5;
      4'b0110 : _zz_PmpPlugin_dGuard_hits_12 = PmpPlugin_mask_6;
      4'b0111 : _zz_PmpPlugin_dGuard_hits_12 = PmpPlugin_mask_7;
      4'b1000 : _zz_PmpPlugin_dGuard_hits_12 = PmpPlugin_mask_8;
      4'b1001 : _zz_PmpPlugin_dGuard_hits_12 = PmpPlugin_mask_9;
      4'b1010 : _zz_PmpPlugin_dGuard_hits_12 = PmpPlugin_mask_10;
      4'b1011 : _zz_PmpPlugin_dGuard_hits_12 = PmpPlugin_mask_11;
      4'b1100 : _zz_PmpPlugin_dGuard_hits_12 = PmpPlugin_mask_12;
      4'b1101 : _zz_PmpPlugin_dGuard_hits_12 = PmpPlugin_mask_13;
      4'b1110 : _zz_PmpPlugin_dGuard_hits_12 = PmpPlugin_mask_14;
      default : _zz_PmpPlugin_dGuard_hits_12 = PmpPlugin_mask_15;
    endcase
  end

  always @(*) begin
    case(_zz_PmpPlugin_dGuard_hits_12_3)
      4'b0000 : _zz_PmpPlugin_dGuard_hits_12_2 = PmpPlugin_base_0;
      4'b0001 : _zz_PmpPlugin_dGuard_hits_12_2 = PmpPlugin_base_1;
      4'b0010 : _zz_PmpPlugin_dGuard_hits_12_2 = PmpPlugin_base_2;
      4'b0011 : _zz_PmpPlugin_dGuard_hits_12_2 = PmpPlugin_base_3;
      4'b0100 : _zz_PmpPlugin_dGuard_hits_12_2 = PmpPlugin_base_4;
      4'b0101 : _zz_PmpPlugin_dGuard_hits_12_2 = PmpPlugin_base_5;
      4'b0110 : _zz_PmpPlugin_dGuard_hits_12_2 = PmpPlugin_base_6;
      4'b0111 : _zz_PmpPlugin_dGuard_hits_12_2 = PmpPlugin_base_7;
      4'b1000 : _zz_PmpPlugin_dGuard_hits_12_2 = PmpPlugin_base_8;
      4'b1001 : _zz_PmpPlugin_dGuard_hits_12_2 = PmpPlugin_base_9;
      4'b1010 : _zz_PmpPlugin_dGuard_hits_12_2 = PmpPlugin_base_10;
      4'b1011 : _zz_PmpPlugin_dGuard_hits_12_2 = PmpPlugin_base_11;
      4'b1100 : _zz_PmpPlugin_dGuard_hits_12_2 = PmpPlugin_base_12;
      4'b1101 : _zz_PmpPlugin_dGuard_hits_12_2 = PmpPlugin_base_13;
      4'b1110 : _zz_PmpPlugin_dGuard_hits_12_2 = PmpPlugin_base_14;
      default : _zz_PmpPlugin_dGuard_hits_12_2 = PmpPlugin_base_15;
    endcase
  end

  always @(*) begin
    case(_zz_PmpPlugin_dGuard_hits_13_1)
      4'b0000 : _zz_PmpPlugin_dGuard_hits_13 = PmpPlugin_mask_0;
      4'b0001 : _zz_PmpPlugin_dGuard_hits_13 = PmpPlugin_mask_1;
      4'b0010 : _zz_PmpPlugin_dGuard_hits_13 = PmpPlugin_mask_2;
      4'b0011 : _zz_PmpPlugin_dGuard_hits_13 = PmpPlugin_mask_3;
      4'b0100 : _zz_PmpPlugin_dGuard_hits_13 = PmpPlugin_mask_4;
      4'b0101 : _zz_PmpPlugin_dGuard_hits_13 = PmpPlugin_mask_5;
      4'b0110 : _zz_PmpPlugin_dGuard_hits_13 = PmpPlugin_mask_6;
      4'b0111 : _zz_PmpPlugin_dGuard_hits_13 = PmpPlugin_mask_7;
      4'b1000 : _zz_PmpPlugin_dGuard_hits_13 = PmpPlugin_mask_8;
      4'b1001 : _zz_PmpPlugin_dGuard_hits_13 = PmpPlugin_mask_9;
      4'b1010 : _zz_PmpPlugin_dGuard_hits_13 = PmpPlugin_mask_10;
      4'b1011 : _zz_PmpPlugin_dGuard_hits_13 = PmpPlugin_mask_11;
      4'b1100 : _zz_PmpPlugin_dGuard_hits_13 = PmpPlugin_mask_12;
      4'b1101 : _zz_PmpPlugin_dGuard_hits_13 = PmpPlugin_mask_13;
      4'b1110 : _zz_PmpPlugin_dGuard_hits_13 = PmpPlugin_mask_14;
      default : _zz_PmpPlugin_dGuard_hits_13 = PmpPlugin_mask_15;
    endcase
  end

  always @(*) begin
    case(_zz_PmpPlugin_dGuard_hits_13_3)
      4'b0000 : _zz_PmpPlugin_dGuard_hits_13_2 = PmpPlugin_base_0;
      4'b0001 : _zz_PmpPlugin_dGuard_hits_13_2 = PmpPlugin_base_1;
      4'b0010 : _zz_PmpPlugin_dGuard_hits_13_2 = PmpPlugin_base_2;
      4'b0011 : _zz_PmpPlugin_dGuard_hits_13_2 = PmpPlugin_base_3;
      4'b0100 : _zz_PmpPlugin_dGuard_hits_13_2 = PmpPlugin_base_4;
      4'b0101 : _zz_PmpPlugin_dGuard_hits_13_2 = PmpPlugin_base_5;
      4'b0110 : _zz_PmpPlugin_dGuard_hits_13_2 = PmpPlugin_base_6;
      4'b0111 : _zz_PmpPlugin_dGuard_hits_13_2 = PmpPlugin_base_7;
      4'b1000 : _zz_PmpPlugin_dGuard_hits_13_2 = PmpPlugin_base_8;
      4'b1001 : _zz_PmpPlugin_dGuard_hits_13_2 = PmpPlugin_base_9;
      4'b1010 : _zz_PmpPlugin_dGuard_hits_13_2 = PmpPlugin_base_10;
      4'b1011 : _zz_PmpPlugin_dGuard_hits_13_2 = PmpPlugin_base_11;
      4'b1100 : _zz_PmpPlugin_dGuard_hits_13_2 = PmpPlugin_base_12;
      4'b1101 : _zz_PmpPlugin_dGuard_hits_13_2 = PmpPlugin_base_13;
      4'b1110 : _zz_PmpPlugin_dGuard_hits_13_2 = PmpPlugin_base_14;
      default : _zz_PmpPlugin_dGuard_hits_13_2 = PmpPlugin_base_15;
    endcase
  end

  always @(*) begin
    case(_zz_PmpPlugin_dGuard_hits_14_1)
      4'b0000 : _zz_PmpPlugin_dGuard_hits_14 = PmpPlugin_mask_0;
      4'b0001 : _zz_PmpPlugin_dGuard_hits_14 = PmpPlugin_mask_1;
      4'b0010 : _zz_PmpPlugin_dGuard_hits_14 = PmpPlugin_mask_2;
      4'b0011 : _zz_PmpPlugin_dGuard_hits_14 = PmpPlugin_mask_3;
      4'b0100 : _zz_PmpPlugin_dGuard_hits_14 = PmpPlugin_mask_4;
      4'b0101 : _zz_PmpPlugin_dGuard_hits_14 = PmpPlugin_mask_5;
      4'b0110 : _zz_PmpPlugin_dGuard_hits_14 = PmpPlugin_mask_6;
      4'b0111 : _zz_PmpPlugin_dGuard_hits_14 = PmpPlugin_mask_7;
      4'b1000 : _zz_PmpPlugin_dGuard_hits_14 = PmpPlugin_mask_8;
      4'b1001 : _zz_PmpPlugin_dGuard_hits_14 = PmpPlugin_mask_9;
      4'b1010 : _zz_PmpPlugin_dGuard_hits_14 = PmpPlugin_mask_10;
      4'b1011 : _zz_PmpPlugin_dGuard_hits_14 = PmpPlugin_mask_11;
      4'b1100 : _zz_PmpPlugin_dGuard_hits_14 = PmpPlugin_mask_12;
      4'b1101 : _zz_PmpPlugin_dGuard_hits_14 = PmpPlugin_mask_13;
      4'b1110 : _zz_PmpPlugin_dGuard_hits_14 = PmpPlugin_mask_14;
      default : _zz_PmpPlugin_dGuard_hits_14 = PmpPlugin_mask_15;
    endcase
  end

  always @(*) begin
    case(_zz_PmpPlugin_dGuard_hits_14_3)
      4'b0000 : _zz_PmpPlugin_dGuard_hits_14_2 = PmpPlugin_base_0;
      4'b0001 : _zz_PmpPlugin_dGuard_hits_14_2 = PmpPlugin_base_1;
      4'b0010 : _zz_PmpPlugin_dGuard_hits_14_2 = PmpPlugin_base_2;
      4'b0011 : _zz_PmpPlugin_dGuard_hits_14_2 = PmpPlugin_base_3;
      4'b0100 : _zz_PmpPlugin_dGuard_hits_14_2 = PmpPlugin_base_4;
      4'b0101 : _zz_PmpPlugin_dGuard_hits_14_2 = PmpPlugin_base_5;
      4'b0110 : _zz_PmpPlugin_dGuard_hits_14_2 = PmpPlugin_base_6;
      4'b0111 : _zz_PmpPlugin_dGuard_hits_14_2 = PmpPlugin_base_7;
      4'b1000 : _zz_PmpPlugin_dGuard_hits_14_2 = PmpPlugin_base_8;
      4'b1001 : _zz_PmpPlugin_dGuard_hits_14_2 = PmpPlugin_base_9;
      4'b1010 : _zz_PmpPlugin_dGuard_hits_14_2 = PmpPlugin_base_10;
      4'b1011 : _zz_PmpPlugin_dGuard_hits_14_2 = PmpPlugin_base_11;
      4'b1100 : _zz_PmpPlugin_dGuard_hits_14_2 = PmpPlugin_base_12;
      4'b1101 : _zz_PmpPlugin_dGuard_hits_14_2 = PmpPlugin_base_13;
      4'b1110 : _zz_PmpPlugin_dGuard_hits_14_2 = PmpPlugin_base_14;
      default : _zz_PmpPlugin_dGuard_hits_14_2 = PmpPlugin_base_15;
    endcase
  end

  always @(*) begin
    case(_zz_PmpPlugin_dGuard_hits_15_1)
      4'b0000 : _zz_PmpPlugin_dGuard_hits_15 = PmpPlugin_mask_0;
      4'b0001 : _zz_PmpPlugin_dGuard_hits_15 = PmpPlugin_mask_1;
      4'b0010 : _zz_PmpPlugin_dGuard_hits_15 = PmpPlugin_mask_2;
      4'b0011 : _zz_PmpPlugin_dGuard_hits_15 = PmpPlugin_mask_3;
      4'b0100 : _zz_PmpPlugin_dGuard_hits_15 = PmpPlugin_mask_4;
      4'b0101 : _zz_PmpPlugin_dGuard_hits_15 = PmpPlugin_mask_5;
      4'b0110 : _zz_PmpPlugin_dGuard_hits_15 = PmpPlugin_mask_6;
      4'b0111 : _zz_PmpPlugin_dGuard_hits_15 = PmpPlugin_mask_7;
      4'b1000 : _zz_PmpPlugin_dGuard_hits_15 = PmpPlugin_mask_8;
      4'b1001 : _zz_PmpPlugin_dGuard_hits_15 = PmpPlugin_mask_9;
      4'b1010 : _zz_PmpPlugin_dGuard_hits_15 = PmpPlugin_mask_10;
      4'b1011 : _zz_PmpPlugin_dGuard_hits_15 = PmpPlugin_mask_11;
      4'b1100 : _zz_PmpPlugin_dGuard_hits_15 = PmpPlugin_mask_12;
      4'b1101 : _zz_PmpPlugin_dGuard_hits_15 = PmpPlugin_mask_13;
      4'b1110 : _zz_PmpPlugin_dGuard_hits_15 = PmpPlugin_mask_14;
      default : _zz_PmpPlugin_dGuard_hits_15 = PmpPlugin_mask_15;
    endcase
  end

  always @(*) begin
    case(_zz_PmpPlugin_dGuard_hits_15_3)
      4'b0000 : _zz_PmpPlugin_dGuard_hits_15_2 = PmpPlugin_base_0;
      4'b0001 : _zz_PmpPlugin_dGuard_hits_15_2 = PmpPlugin_base_1;
      4'b0010 : _zz_PmpPlugin_dGuard_hits_15_2 = PmpPlugin_base_2;
      4'b0011 : _zz_PmpPlugin_dGuard_hits_15_2 = PmpPlugin_base_3;
      4'b0100 : _zz_PmpPlugin_dGuard_hits_15_2 = PmpPlugin_base_4;
      4'b0101 : _zz_PmpPlugin_dGuard_hits_15_2 = PmpPlugin_base_5;
      4'b0110 : _zz_PmpPlugin_dGuard_hits_15_2 = PmpPlugin_base_6;
      4'b0111 : _zz_PmpPlugin_dGuard_hits_15_2 = PmpPlugin_base_7;
      4'b1000 : _zz_PmpPlugin_dGuard_hits_15_2 = PmpPlugin_base_8;
      4'b1001 : _zz_PmpPlugin_dGuard_hits_15_2 = PmpPlugin_base_9;
      4'b1010 : _zz_PmpPlugin_dGuard_hits_15_2 = PmpPlugin_base_10;
      4'b1011 : _zz_PmpPlugin_dGuard_hits_15_2 = PmpPlugin_base_11;
      4'b1100 : _zz_PmpPlugin_dGuard_hits_15_2 = PmpPlugin_base_12;
      4'b1101 : _zz_PmpPlugin_dGuard_hits_15_2 = PmpPlugin_base_13;
      4'b1110 : _zz_PmpPlugin_dGuard_hits_15_2 = PmpPlugin_base_14;
      default : _zz_PmpPlugin_dGuard_hits_15_2 = PmpPlugin_base_15;
    endcase
  end

  always @(*) begin
    case(_zz_DBusCachedPlugin_mmuBus_rsp_allowRead_18)
      4'b0000 : _zz_DBusCachedPlugin_mmuBus_rsp_allowRead_17 = PmpPlugin_pmpcfg_0[0];
      4'b0001 : _zz_DBusCachedPlugin_mmuBus_rsp_allowRead_17 = PmpPlugin_pmpcfg_1[0];
      4'b0010 : _zz_DBusCachedPlugin_mmuBus_rsp_allowRead_17 = PmpPlugin_pmpcfg_2[0];
      4'b0011 : _zz_DBusCachedPlugin_mmuBus_rsp_allowRead_17 = PmpPlugin_pmpcfg_3[0];
      4'b0100 : _zz_DBusCachedPlugin_mmuBus_rsp_allowRead_17 = PmpPlugin_pmpcfg_4[0];
      4'b0101 : _zz_DBusCachedPlugin_mmuBus_rsp_allowRead_17 = PmpPlugin_pmpcfg_5[0];
      4'b0110 : _zz_DBusCachedPlugin_mmuBus_rsp_allowRead_17 = PmpPlugin_pmpcfg_6[0];
      4'b0111 : _zz_DBusCachedPlugin_mmuBus_rsp_allowRead_17 = PmpPlugin_pmpcfg_7[0];
      4'b1000 : _zz_DBusCachedPlugin_mmuBus_rsp_allowRead_17 = PmpPlugin_pmpcfg_8[0];
      4'b1001 : _zz_DBusCachedPlugin_mmuBus_rsp_allowRead_17 = PmpPlugin_pmpcfg_9[0];
      4'b1010 : _zz_DBusCachedPlugin_mmuBus_rsp_allowRead_17 = PmpPlugin_pmpcfg_10[0];
      4'b1011 : _zz_DBusCachedPlugin_mmuBus_rsp_allowRead_17 = PmpPlugin_pmpcfg_11[0];
      4'b1100 : _zz_DBusCachedPlugin_mmuBus_rsp_allowRead_17 = PmpPlugin_pmpcfg_12[0];
      4'b1101 : _zz_DBusCachedPlugin_mmuBus_rsp_allowRead_17 = PmpPlugin_pmpcfg_13[0];
      4'b1110 : _zz_DBusCachedPlugin_mmuBus_rsp_allowRead_17 = PmpPlugin_pmpcfg_14[0];
      default : _zz_DBusCachedPlugin_mmuBus_rsp_allowRead_17 = PmpPlugin_pmpcfg_15[0];
    endcase
  end

  always @(*) begin
    case(_zz_DBusCachedPlugin_mmuBus_rsp_allowWrite_18)
      4'b0000 : _zz_DBusCachedPlugin_mmuBus_rsp_allowWrite_17 = PmpPlugin_pmpcfg_0[1];
      4'b0001 : _zz_DBusCachedPlugin_mmuBus_rsp_allowWrite_17 = PmpPlugin_pmpcfg_1[1];
      4'b0010 : _zz_DBusCachedPlugin_mmuBus_rsp_allowWrite_17 = PmpPlugin_pmpcfg_2[1];
      4'b0011 : _zz_DBusCachedPlugin_mmuBus_rsp_allowWrite_17 = PmpPlugin_pmpcfg_3[1];
      4'b0100 : _zz_DBusCachedPlugin_mmuBus_rsp_allowWrite_17 = PmpPlugin_pmpcfg_4[1];
      4'b0101 : _zz_DBusCachedPlugin_mmuBus_rsp_allowWrite_17 = PmpPlugin_pmpcfg_5[1];
      4'b0110 : _zz_DBusCachedPlugin_mmuBus_rsp_allowWrite_17 = PmpPlugin_pmpcfg_6[1];
      4'b0111 : _zz_DBusCachedPlugin_mmuBus_rsp_allowWrite_17 = PmpPlugin_pmpcfg_7[1];
      4'b1000 : _zz_DBusCachedPlugin_mmuBus_rsp_allowWrite_17 = PmpPlugin_pmpcfg_8[1];
      4'b1001 : _zz_DBusCachedPlugin_mmuBus_rsp_allowWrite_17 = PmpPlugin_pmpcfg_9[1];
      4'b1010 : _zz_DBusCachedPlugin_mmuBus_rsp_allowWrite_17 = PmpPlugin_pmpcfg_10[1];
      4'b1011 : _zz_DBusCachedPlugin_mmuBus_rsp_allowWrite_17 = PmpPlugin_pmpcfg_11[1];
      4'b1100 : _zz_DBusCachedPlugin_mmuBus_rsp_allowWrite_17 = PmpPlugin_pmpcfg_12[1];
      4'b1101 : _zz_DBusCachedPlugin_mmuBus_rsp_allowWrite_17 = PmpPlugin_pmpcfg_13[1];
      4'b1110 : _zz_DBusCachedPlugin_mmuBus_rsp_allowWrite_17 = PmpPlugin_pmpcfg_14[1];
      default : _zz_DBusCachedPlugin_mmuBus_rsp_allowWrite_17 = PmpPlugin_pmpcfg_15[1];
    endcase
  end

  always @(*) begin
    case(_zz_PmpPlugin_iGuard_hits_0_2)
      4'b0000 : _zz_PmpPlugin_iGuard_hits_0_1 = PmpPlugin_mask_0;
      4'b0001 : _zz_PmpPlugin_iGuard_hits_0_1 = PmpPlugin_mask_1;
      4'b0010 : _zz_PmpPlugin_iGuard_hits_0_1 = PmpPlugin_mask_2;
      4'b0011 : _zz_PmpPlugin_iGuard_hits_0_1 = PmpPlugin_mask_3;
      4'b0100 : _zz_PmpPlugin_iGuard_hits_0_1 = PmpPlugin_mask_4;
      4'b0101 : _zz_PmpPlugin_iGuard_hits_0_1 = PmpPlugin_mask_5;
      4'b0110 : _zz_PmpPlugin_iGuard_hits_0_1 = PmpPlugin_mask_6;
      4'b0111 : _zz_PmpPlugin_iGuard_hits_0_1 = PmpPlugin_mask_7;
      4'b1000 : _zz_PmpPlugin_iGuard_hits_0_1 = PmpPlugin_mask_8;
      4'b1001 : _zz_PmpPlugin_iGuard_hits_0_1 = PmpPlugin_mask_9;
      4'b1010 : _zz_PmpPlugin_iGuard_hits_0_1 = PmpPlugin_mask_10;
      4'b1011 : _zz_PmpPlugin_iGuard_hits_0_1 = PmpPlugin_mask_11;
      4'b1100 : _zz_PmpPlugin_iGuard_hits_0_1 = PmpPlugin_mask_12;
      4'b1101 : _zz_PmpPlugin_iGuard_hits_0_1 = PmpPlugin_mask_13;
      4'b1110 : _zz_PmpPlugin_iGuard_hits_0_1 = PmpPlugin_mask_14;
      default : _zz_PmpPlugin_iGuard_hits_0_1 = PmpPlugin_mask_15;
    endcase
  end

  always @(*) begin
    case(_zz_PmpPlugin_iGuard_hits_0_4)
      4'b0000 : _zz_PmpPlugin_iGuard_hits_0_3 = PmpPlugin_base_0;
      4'b0001 : _zz_PmpPlugin_iGuard_hits_0_3 = PmpPlugin_base_1;
      4'b0010 : _zz_PmpPlugin_iGuard_hits_0_3 = PmpPlugin_base_2;
      4'b0011 : _zz_PmpPlugin_iGuard_hits_0_3 = PmpPlugin_base_3;
      4'b0100 : _zz_PmpPlugin_iGuard_hits_0_3 = PmpPlugin_base_4;
      4'b0101 : _zz_PmpPlugin_iGuard_hits_0_3 = PmpPlugin_base_5;
      4'b0110 : _zz_PmpPlugin_iGuard_hits_0_3 = PmpPlugin_base_6;
      4'b0111 : _zz_PmpPlugin_iGuard_hits_0_3 = PmpPlugin_base_7;
      4'b1000 : _zz_PmpPlugin_iGuard_hits_0_3 = PmpPlugin_base_8;
      4'b1001 : _zz_PmpPlugin_iGuard_hits_0_3 = PmpPlugin_base_9;
      4'b1010 : _zz_PmpPlugin_iGuard_hits_0_3 = PmpPlugin_base_10;
      4'b1011 : _zz_PmpPlugin_iGuard_hits_0_3 = PmpPlugin_base_11;
      4'b1100 : _zz_PmpPlugin_iGuard_hits_0_3 = PmpPlugin_base_12;
      4'b1101 : _zz_PmpPlugin_iGuard_hits_0_3 = PmpPlugin_base_13;
      4'b1110 : _zz_PmpPlugin_iGuard_hits_0_3 = PmpPlugin_base_14;
      default : _zz_PmpPlugin_iGuard_hits_0_3 = PmpPlugin_base_15;
    endcase
  end

  always @(*) begin
    case(_zz_PmpPlugin_iGuard_hits_1_1)
      4'b0000 : _zz_PmpPlugin_iGuard_hits_1 = PmpPlugin_mask_0;
      4'b0001 : _zz_PmpPlugin_iGuard_hits_1 = PmpPlugin_mask_1;
      4'b0010 : _zz_PmpPlugin_iGuard_hits_1 = PmpPlugin_mask_2;
      4'b0011 : _zz_PmpPlugin_iGuard_hits_1 = PmpPlugin_mask_3;
      4'b0100 : _zz_PmpPlugin_iGuard_hits_1 = PmpPlugin_mask_4;
      4'b0101 : _zz_PmpPlugin_iGuard_hits_1 = PmpPlugin_mask_5;
      4'b0110 : _zz_PmpPlugin_iGuard_hits_1 = PmpPlugin_mask_6;
      4'b0111 : _zz_PmpPlugin_iGuard_hits_1 = PmpPlugin_mask_7;
      4'b1000 : _zz_PmpPlugin_iGuard_hits_1 = PmpPlugin_mask_8;
      4'b1001 : _zz_PmpPlugin_iGuard_hits_1 = PmpPlugin_mask_9;
      4'b1010 : _zz_PmpPlugin_iGuard_hits_1 = PmpPlugin_mask_10;
      4'b1011 : _zz_PmpPlugin_iGuard_hits_1 = PmpPlugin_mask_11;
      4'b1100 : _zz_PmpPlugin_iGuard_hits_1 = PmpPlugin_mask_12;
      4'b1101 : _zz_PmpPlugin_iGuard_hits_1 = PmpPlugin_mask_13;
      4'b1110 : _zz_PmpPlugin_iGuard_hits_1 = PmpPlugin_mask_14;
      default : _zz_PmpPlugin_iGuard_hits_1 = PmpPlugin_mask_15;
    endcase
  end

  always @(*) begin
    case(_zz_PmpPlugin_iGuard_hits_1_3)
      4'b0000 : _zz_PmpPlugin_iGuard_hits_1_2 = PmpPlugin_base_0;
      4'b0001 : _zz_PmpPlugin_iGuard_hits_1_2 = PmpPlugin_base_1;
      4'b0010 : _zz_PmpPlugin_iGuard_hits_1_2 = PmpPlugin_base_2;
      4'b0011 : _zz_PmpPlugin_iGuard_hits_1_2 = PmpPlugin_base_3;
      4'b0100 : _zz_PmpPlugin_iGuard_hits_1_2 = PmpPlugin_base_4;
      4'b0101 : _zz_PmpPlugin_iGuard_hits_1_2 = PmpPlugin_base_5;
      4'b0110 : _zz_PmpPlugin_iGuard_hits_1_2 = PmpPlugin_base_6;
      4'b0111 : _zz_PmpPlugin_iGuard_hits_1_2 = PmpPlugin_base_7;
      4'b1000 : _zz_PmpPlugin_iGuard_hits_1_2 = PmpPlugin_base_8;
      4'b1001 : _zz_PmpPlugin_iGuard_hits_1_2 = PmpPlugin_base_9;
      4'b1010 : _zz_PmpPlugin_iGuard_hits_1_2 = PmpPlugin_base_10;
      4'b1011 : _zz_PmpPlugin_iGuard_hits_1_2 = PmpPlugin_base_11;
      4'b1100 : _zz_PmpPlugin_iGuard_hits_1_2 = PmpPlugin_base_12;
      4'b1101 : _zz_PmpPlugin_iGuard_hits_1_2 = PmpPlugin_base_13;
      4'b1110 : _zz_PmpPlugin_iGuard_hits_1_2 = PmpPlugin_base_14;
      default : _zz_PmpPlugin_iGuard_hits_1_2 = PmpPlugin_base_15;
    endcase
  end

  always @(*) begin
    case(_zz_PmpPlugin_iGuard_hits_2_1)
      4'b0000 : _zz_PmpPlugin_iGuard_hits_2 = PmpPlugin_mask_0;
      4'b0001 : _zz_PmpPlugin_iGuard_hits_2 = PmpPlugin_mask_1;
      4'b0010 : _zz_PmpPlugin_iGuard_hits_2 = PmpPlugin_mask_2;
      4'b0011 : _zz_PmpPlugin_iGuard_hits_2 = PmpPlugin_mask_3;
      4'b0100 : _zz_PmpPlugin_iGuard_hits_2 = PmpPlugin_mask_4;
      4'b0101 : _zz_PmpPlugin_iGuard_hits_2 = PmpPlugin_mask_5;
      4'b0110 : _zz_PmpPlugin_iGuard_hits_2 = PmpPlugin_mask_6;
      4'b0111 : _zz_PmpPlugin_iGuard_hits_2 = PmpPlugin_mask_7;
      4'b1000 : _zz_PmpPlugin_iGuard_hits_2 = PmpPlugin_mask_8;
      4'b1001 : _zz_PmpPlugin_iGuard_hits_2 = PmpPlugin_mask_9;
      4'b1010 : _zz_PmpPlugin_iGuard_hits_2 = PmpPlugin_mask_10;
      4'b1011 : _zz_PmpPlugin_iGuard_hits_2 = PmpPlugin_mask_11;
      4'b1100 : _zz_PmpPlugin_iGuard_hits_2 = PmpPlugin_mask_12;
      4'b1101 : _zz_PmpPlugin_iGuard_hits_2 = PmpPlugin_mask_13;
      4'b1110 : _zz_PmpPlugin_iGuard_hits_2 = PmpPlugin_mask_14;
      default : _zz_PmpPlugin_iGuard_hits_2 = PmpPlugin_mask_15;
    endcase
  end

  always @(*) begin
    case(_zz_PmpPlugin_iGuard_hits_2_3)
      4'b0000 : _zz_PmpPlugin_iGuard_hits_2_2 = PmpPlugin_base_0;
      4'b0001 : _zz_PmpPlugin_iGuard_hits_2_2 = PmpPlugin_base_1;
      4'b0010 : _zz_PmpPlugin_iGuard_hits_2_2 = PmpPlugin_base_2;
      4'b0011 : _zz_PmpPlugin_iGuard_hits_2_2 = PmpPlugin_base_3;
      4'b0100 : _zz_PmpPlugin_iGuard_hits_2_2 = PmpPlugin_base_4;
      4'b0101 : _zz_PmpPlugin_iGuard_hits_2_2 = PmpPlugin_base_5;
      4'b0110 : _zz_PmpPlugin_iGuard_hits_2_2 = PmpPlugin_base_6;
      4'b0111 : _zz_PmpPlugin_iGuard_hits_2_2 = PmpPlugin_base_7;
      4'b1000 : _zz_PmpPlugin_iGuard_hits_2_2 = PmpPlugin_base_8;
      4'b1001 : _zz_PmpPlugin_iGuard_hits_2_2 = PmpPlugin_base_9;
      4'b1010 : _zz_PmpPlugin_iGuard_hits_2_2 = PmpPlugin_base_10;
      4'b1011 : _zz_PmpPlugin_iGuard_hits_2_2 = PmpPlugin_base_11;
      4'b1100 : _zz_PmpPlugin_iGuard_hits_2_2 = PmpPlugin_base_12;
      4'b1101 : _zz_PmpPlugin_iGuard_hits_2_2 = PmpPlugin_base_13;
      4'b1110 : _zz_PmpPlugin_iGuard_hits_2_2 = PmpPlugin_base_14;
      default : _zz_PmpPlugin_iGuard_hits_2_2 = PmpPlugin_base_15;
    endcase
  end

  always @(*) begin
    case(_zz_PmpPlugin_iGuard_hits_3_1)
      4'b0000 : _zz_PmpPlugin_iGuard_hits_3 = PmpPlugin_mask_0;
      4'b0001 : _zz_PmpPlugin_iGuard_hits_3 = PmpPlugin_mask_1;
      4'b0010 : _zz_PmpPlugin_iGuard_hits_3 = PmpPlugin_mask_2;
      4'b0011 : _zz_PmpPlugin_iGuard_hits_3 = PmpPlugin_mask_3;
      4'b0100 : _zz_PmpPlugin_iGuard_hits_3 = PmpPlugin_mask_4;
      4'b0101 : _zz_PmpPlugin_iGuard_hits_3 = PmpPlugin_mask_5;
      4'b0110 : _zz_PmpPlugin_iGuard_hits_3 = PmpPlugin_mask_6;
      4'b0111 : _zz_PmpPlugin_iGuard_hits_3 = PmpPlugin_mask_7;
      4'b1000 : _zz_PmpPlugin_iGuard_hits_3 = PmpPlugin_mask_8;
      4'b1001 : _zz_PmpPlugin_iGuard_hits_3 = PmpPlugin_mask_9;
      4'b1010 : _zz_PmpPlugin_iGuard_hits_3 = PmpPlugin_mask_10;
      4'b1011 : _zz_PmpPlugin_iGuard_hits_3 = PmpPlugin_mask_11;
      4'b1100 : _zz_PmpPlugin_iGuard_hits_3 = PmpPlugin_mask_12;
      4'b1101 : _zz_PmpPlugin_iGuard_hits_3 = PmpPlugin_mask_13;
      4'b1110 : _zz_PmpPlugin_iGuard_hits_3 = PmpPlugin_mask_14;
      default : _zz_PmpPlugin_iGuard_hits_3 = PmpPlugin_mask_15;
    endcase
  end

  always @(*) begin
    case(_zz_PmpPlugin_iGuard_hits_3_3)
      4'b0000 : _zz_PmpPlugin_iGuard_hits_3_2 = PmpPlugin_base_0;
      4'b0001 : _zz_PmpPlugin_iGuard_hits_3_2 = PmpPlugin_base_1;
      4'b0010 : _zz_PmpPlugin_iGuard_hits_3_2 = PmpPlugin_base_2;
      4'b0011 : _zz_PmpPlugin_iGuard_hits_3_2 = PmpPlugin_base_3;
      4'b0100 : _zz_PmpPlugin_iGuard_hits_3_2 = PmpPlugin_base_4;
      4'b0101 : _zz_PmpPlugin_iGuard_hits_3_2 = PmpPlugin_base_5;
      4'b0110 : _zz_PmpPlugin_iGuard_hits_3_2 = PmpPlugin_base_6;
      4'b0111 : _zz_PmpPlugin_iGuard_hits_3_2 = PmpPlugin_base_7;
      4'b1000 : _zz_PmpPlugin_iGuard_hits_3_2 = PmpPlugin_base_8;
      4'b1001 : _zz_PmpPlugin_iGuard_hits_3_2 = PmpPlugin_base_9;
      4'b1010 : _zz_PmpPlugin_iGuard_hits_3_2 = PmpPlugin_base_10;
      4'b1011 : _zz_PmpPlugin_iGuard_hits_3_2 = PmpPlugin_base_11;
      4'b1100 : _zz_PmpPlugin_iGuard_hits_3_2 = PmpPlugin_base_12;
      4'b1101 : _zz_PmpPlugin_iGuard_hits_3_2 = PmpPlugin_base_13;
      4'b1110 : _zz_PmpPlugin_iGuard_hits_3_2 = PmpPlugin_base_14;
      default : _zz_PmpPlugin_iGuard_hits_3_2 = PmpPlugin_base_15;
    endcase
  end

  always @(*) begin
    case(_zz_PmpPlugin_iGuard_hits_4_1)
      4'b0000 : _zz_PmpPlugin_iGuard_hits_4 = PmpPlugin_mask_0;
      4'b0001 : _zz_PmpPlugin_iGuard_hits_4 = PmpPlugin_mask_1;
      4'b0010 : _zz_PmpPlugin_iGuard_hits_4 = PmpPlugin_mask_2;
      4'b0011 : _zz_PmpPlugin_iGuard_hits_4 = PmpPlugin_mask_3;
      4'b0100 : _zz_PmpPlugin_iGuard_hits_4 = PmpPlugin_mask_4;
      4'b0101 : _zz_PmpPlugin_iGuard_hits_4 = PmpPlugin_mask_5;
      4'b0110 : _zz_PmpPlugin_iGuard_hits_4 = PmpPlugin_mask_6;
      4'b0111 : _zz_PmpPlugin_iGuard_hits_4 = PmpPlugin_mask_7;
      4'b1000 : _zz_PmpPlugin_iGuard_hits_4 = PmpPlugin_mask_8;
      4'b1001 : _zz_PmpPlugin_iGuard_hits_4 = PmpPlugin_mask_9;
      4'b1010 : _zz_PmpPlugin_iGuard_hits_4 = PmpPlugin_mask_10;
      4'b1011 : _zz_PmpPlugin_iGuard_hits_4 = PmpPlugin_mask_11;
      4'b1100 : _zz_PmpPlugin_iGuard_hits_4 = PmpPlugin_mask_12;
      4'b1101 : _zz_PmpPlugin_iGuard_hits_4 = PmpPlugin_mask_13;
      4'b1110 : _zz_PmpPlugin_iGuard_hits_4 = PmpPlugin_mask_14;
      default : _zz_PmpPlugin_iGuard_hits_4 = PmpPlugin_mask_15;
    endcase
  end

  always @(*) begin
    case(_zz_PmpPlugin_iGuard_hits_4_3)
      4'b0000 : _zz_PmpPlugin_iGuard_hits_4_2 = PmpPlugin_base_0;
      4'b0001 : _zz_PmpPlugin_iGuard_hits_4_2 = PmpPlugin_base_1;
      4'b0010 : _zz_PmpPlugin_iGuard_hits_4_2 = PmpPlugin_base_2;
      4'b0011 : _zz_PmpPlugin_iGuard_hits_4_2 = PmpPlugin_base_3;
      4'b0100 : _zz_PmpPlugin_iGuard_hits_4_2 = PmpPlugin_base_4;
      4'b0101 : _zz_PmpPlugin_iGuard_hits_4_2 = PmpPlugin_base_5;
      4'b0110 : _zz_PmpPlugin_iGuard_hits_4_2 = PmpPlugin_base_6;
      4'b0111 : _zz_PmpPlugin_iGuard_hits_4_2 = PmpPlugin_base_7;
      4'b1000 : _zz_PmpPlugin_iGuard_hits_4_2 = PmpPlugin_base_8;
      4'b1001 : _zz_PmpPlugin_iGuard_hits_4_2 = PmpPlugin_base_9;
      4'b1010 : _zz_PmpPlugin_iGuard_hits_4_2 = PmpPlugin_base_10;
      4'b1011 : _zz_PmpPlugin_iGuard_hits_4_2 = PmpPlugin_base_11;
      4'b1100 : _zz_PmpPlugin_iGuard_hits_4_2 = PmpPlugin_base_12;
      4'b1101 : _zz_PmpPlugin_iGuard_hits_4_2 = PmpPlugin_base_13;
      4'b1110 : _zz_PmpPlugin_iGuard_hits_4_2 = PmpPlugin_base_14;
      default : _zz_PmpPlugin_iGuard_hits_4_2 = PmpPlugin_base_15;
    endcase
  end

  always @(*) begin
    case(_zz_PmpPlugin_iGuard_hits_5_1)
      4'b0000 : _zz_PmpPlugin_iGuard_hits_5 = PmpPlugin_mask_0;
      4'b0001 : _zz_PmpPlugin_iGuard_hits_5 = PmpPlugin_mask_1;
      4'b0010 : _zz_PmpPlugin_iGuard_hits_5 = PmpPlugin_mask_2;
      4'b0011 : _zz_PmpPlugin_iGuard_hits_5 = PmpPlugin_mask_3;
      4'b0100 : _zz_PmpPlugin_iGuard_hits_5 = PmpPlugin_mask_4;
      4'b0101 : _zz_PmpPlugin_iGuard_hits_5 = PmpPlugin_mask_5;
      4'b0110 : _zz_PmpPlugin_iGuard_hits_5 = PmpPlugin_mask_6;
      4'b0111 : _zz_PmpPlugin_iGuard_hits_5 = PmpPlugin_mask_7;
      4'b1000 : _zz_PmpPlugin_iGuard_hits_5 = PmpPlugin_mask_8;
      4'b1001 : _zz_PmpPlugin_iGuard_hits_5 = PmpPlugin_mask_9;
      4'b1010 : _zz_PmpPlugin_iGuard_hits_5 = PmpPlugin_mask_10;
      4'b1011 : _zz_PmpPlugin_iGuard_hits_5 = PmpPlugin_mask_11;
      4'b1100 : _zz_PmpPlugin_iGuard_hits_5 = PmpPlugin_mask_12;
      4'b1101 : _zz_PmpPlugin_iGuard_hits_5 = PmpPlugin_mask_13;
      4'b1110 : _zz_PmpPlugin_iGuard_hits_5 = PmpPlugin_mask_14;
      default : _zz_PmpPlugin_iGuard_hits_5 = PmpPlugin_mask_15;
    endcase
  end

  always @(*) begin
    case(_zz_PmpPlugin_iGuard_hits_5_3)
      4'b0000 : _zz_PmpPlugin_iGuard_hits_5_2 = PmpPlugin_base_0;
      4'b0001 : _zz_PmpPlugin_iGuard_hits_5_2 = PmpPlugin_base_1;
      4'b0010 : _zz_PmpPlugin_iGuard_hits_5_2 = PmpPlugin_base_2;
      4'b0011 : _zz_PmpPlugin_iGuard_hits_5_2 = PmpPlugin_base_3;
      4'b0100 : _zz_PmpPlugin_iGuard_hits_5_2 = PmpPlugin_base_4;
      4'b0101 : _zz_PmpPlugin_iGuard_hits_5_2 = PmpPlugin_base_5;
      4'b0110 : _zz_PmpPlugin_iGuard_hits_5_2 = PmpPlugin_base_6;
      4'b0111 : _zz_PmpPlugin_iGuard_hits_5_2 = PmpPlugin_base_7;
      4'b1000 : _zz_PmpPlugin_iGuard_hits_5_2 = PmpPlugin_base_8;
      4'b1001 : _zz_PmpPlugin_iGuard_hits_5_2 = PmpPlugin_base_9;
      4'b1010 : _zz_PmpPlugin_iGuard_hits_5_2 = PmpPlugin_base_10;
      4'b1011 : _zz_PmpPlugin_iGuard_hits_5_2 = PmpPlugin_base_11;
      4'b1100 : _zz_PmpPlugin_iGuard_hits_5_2 = PmpPlugin_base_12;
      4'b1101 : _zz_PmpPlugin_iGuard_hits_5_2 = PmpPlugin_base_13;
      4'b1110 : _zz_PmpPlugin_iGuard_hits_5_2 = PmpPlugin_base_14;
      default : _zz_PmpPlugin_iGuard_hits_5_2 = PmpPlugin_base_15;
    endcase
  end

  always @(*) begin
    case(_zz_PmpPlugin_iGuard_hits_6_1)
      4'b0000 : _zz_PmpPlugin_iGuard_hits_6 = PmpPlugin_mask_0;
      4'b0001 : _zz_PmpPlugin_iGuard_hits_6 = PmpPlugin_mask_1;
      4'b0010 : _zz_PmpPlugin_iGuard_hits_6 = PmpPlugin_mask_2;
      4'b0011 : _zz_PmpPlugin_iGuard_hits_6 = PmpPlugin_mask_3;
      4'b0100 : _zz_PmpPlugin_iGuard_hits_6 = PmpPlugin_mask_4;
      4'b0101 : _zz_PmpPlugin_iGuard_hits_6 = PmpPlugin_mask_5;
      4'b0110 : _zz_PmpPlugin_iGuard_hits_6 = PmpPlugin_mask_6;
      4'b0111 : _zz_PmpPlugin_iGuard_hits_6 = PmpPlugin_mask_7;
      4'b1000 : _zz_PmpPlugin_iGuard_hits_6 = PmpPlugin_mask_8;
      4'b1001 : _zz_PmpPlugin_iGuard_hits_6 = PmpPlugin_mask_9;
      4'b1010 : _zz_PmpPlugin_iGuard_hits_6 = PmpPlugin_mask_10;
      4'b1011 : _zz_PmpPlugin_iGuard_hits_6 = PmpPlugin_mask_11;
      4'b1100 : _zz_PmpPlugin_iGuard_hits_6 = PmpPlugin_mask_12;
      4'b1101 : _zz_PmpPlugin_iGuard_hits_6 = PmpPlugin_mask_13;
      4'b1110 : _zz_PmpPlugin_iGuard_hits_6 = PmpPlugin_mask_14;
      default : _zz_PmpPlugin_iGuard_hits_6 = PmpPlugin_mask_15;
    endcase
  end

  always @(*) begin
    case(_zz_PmpPlugin_iGuard_hits_6_3)
      4'b0000 : _zz_PmpPlugin_iGuard_hits_6_2 = PmpPlugin_base_0;
      4'b0001 : _zz_PmpPlugin_iGuard_hits_6_2 = PmpPlugin_base_1;
      4'b0010 : _zz_PmpPlugin_iGuard_hits_6_2 = PmpPlugin_base_2;
      4'b0011 : _zz_PmpPlugin_iGuard_hits_6_2 = PmpPlugin_base_3;
      4'b0100 : _zz_PmpPlugin_iGuard_hits_6_2 = PmpPlugin_base_4;
      4'b0101 : _zz_PmpPlugin_iGuard_hits_6_2 = PmpPlugin_base_5;
      4'b0110 : _zz_PmpPlugin_iGuard_hits_6_2 = PmpPlugin_base_6;
      4'b0111 : _zz_PmpPlugin_iGuard_hits_6_2 = PmpPlugin_base_7;
      4'b1000 : _zz_PmpPlugin_iGuard_hits_6_2 = PmpPlugin_base_8;
      4'b1001 : _zz_PmpPlugin_iGuard_hits_6_2 = PmpPlugin_base_9;
      4'b1010 : _zz_PmpPlugin_iGuard_hits_6_2 = PmpPlugin_base_10;
      4'b1011 : _zz_PmpPlugin_iGuard_hits_6_2 = PmpPlugin_base_11;
      4'b1100 : _zz_PmpPlugin_iGuard_hits_6_2 = PmpPlugin_base_12;
      4'b1101 : _zz_PmpPlugin_iGuard_hits_6_2 = PmpPlugin_base_13;
      4'b1110 : _zz_PmpPlugin_iGuard_hits_6_2 = PmpPlugin_base_14;
      default : _zz_PmpPlugin_iGuard_hits_6_2 = PmpPlugin_base_15;
    endcase
  end

  always @(*) begin
    case(_zz_PmpPlugin_iGuard_hits_7_1)
      4'b0000 : _zz_PmpPlugin_iGuard_hits_7 = PmpPlugin_mask_0;
      4'b0001 : _zz_PmpPlugin_iGuard_hits_7 = PmpPlugin_mask_1;
      4'b0010 : _zz_PmpPlugin_iGuard_hits_7 = PmpPlugin_mask_2;
      4'b0011 : _zz_PmpPlugin_iGuard_hits_7 = PmpPlugin_mask_3;
      4'b0100 : _zz_PmpPlugin_iGuard_hits_7 = PmpPlugin_mask_4;
      4'b0101 : _zz_PmpPlugin_iGuard_hits_7 = PmpPlugin_mask_5;
      4'b0110 : _zz_PmpPlugin_iGuard_hits_7 = PmpPlugin_mask_6;
      4'b0111 : _zz_PmpPlugin_iGuard_hits_7 = PmpPlugin_mask_7;
      4'b1000 : _zz_PmpPlugin_iGuard_hits_7 = PmpPlugin_mask_8;
      4'b1001 : _zz_PmpPlugin_iGuard_hits_7 = PmpPlugin_mask_9;
      4'b1010 : _zz_PmpPlugin_iGuard_hits_7 = PmpPlugin_mask_10;
      4'b1011 : _zz_PmpPlugin_iGuard_hits_7 = PmpPlugin_mask_11;
      4'b1100 : _zz_PmpPlugin_iGuard_hits_7 = PmpPlugin_mask_12;
      4'b1101 : _zz_PmpPlugin_iGuard_hits_7 = PmpPlugin_mask_13;
      4'b1110 : _zz_PmpPlugin_iGuard_hits_7 = PmpPlugin_mask_14;
      default : _zz_PmpPlugin_iGuard_hits_7 = PmpPlugin_mask_15;
    endcase
  end

  always @(*) begin
    case(_zz_PmpPlugin_iGuard_hits_7_3)
      4'b0000 : _zz_PmpPlugin_iGuard_hits_7_2 = PmpPlugin_base_0;
      4'b0001 : _zz_PmpPlugin_iGuard_hits_7_2 = PmpPlugin_base_1;
      4'b0010 : _zz_PmpPlugin_iGuard_hits_7_2 = PmpPlugin_base_2;
      4'b0011 : _zz_PmpPlugin_iGuard_hits_7_2 = PmpPlugin_base_3;
      4'b0100 : _zz_PmpPlugin_iGuard_hits_7_2 = PmpPlugin_base_4;
      4'b0101 : _zz_PmpPlugin_iGuard_hits_7_2 = PmpPlugin_base_5;
      4'b0110 : _zz_PmpPlugin_iGuard_hits_7_2 = PmpPlugin_base_6;
      4'b0111 : _zz_PmpPlugin_iGuard_hits_7_2 = PmpPlugin_base_7;
      4'b1000 : _zz_PmpPlugin_iGuard_hits_7_2 = PmpPlugin_base_8;
      4'b1001 : _zz_PmpPlugin_iGuard_hits_7_2 = PmpPlugin_base_9;
      4'b1010 : _zz_PmpPlugin_iGuard_hits_7_2 = PmpPlugin_base_10;
      4'b1011 : _zz_PmpPlugin_iGuard_hits_7_2 = PmpPlugin_base_11;
      4'b1100 : _zz_PmpPlugin_iGuard_hits_7_2 = PmpPlugin_base_12;
      4'b1101 : _zz_PmpPlugin_iGuard_hits_7_2 = PmpPlugin_base_13;
      4'b1110 : _zz_PmpPlugin_iGuard_hits_7_2 = PmpPlugin_base_14;
      default : _zz_PmpPlugin_iGuard_hits_7_2 = PmpPlugin_base_15;
    endcase
  end

  always @(*) begin
    case(_zz_PmpPlugin_iGuard_hits_8_1)
      4'b0000 : _zz_PmpPlugin_iGuard_hits_8 = PmpPlugin_mask_0;
      4'b0001 : _zz_PmpPlugin_iGuard_hits_8 = PmpPlugin_mask_1;
      4'b0010 : _zz_PmpPlugin_iGuard_hits_8 = PmpPlugin_mask_2;
      4'b0011 : _zz_PmpPlugin_iGuard_hits_8 = PmpPlugin_mask_3;
      4'b0100 : _zz_PmpPlugin_iGuard_hits_8 = PmpPlugin_mask_4;
      4'b0101 : _zz_PmpPlugin_iGuard_hits_8 = PmpPlugin_mask_5;
      4'b0110 : _zz_PmpPlugin_iGuard_hits_8 = PmpPlugin_mask_6;
      4'b0111 : _zz_PmpPlugin_iGuard_hits_8 = PmpPlugin_mask_7;
      4'b1000 : _zz_PmpPlugin_iGuard_hits_8 = PmpPlugin_mask_8;
      4'b1001 : _zz_PmpPlugin_iGuard_hits_8 = PmpPlugin_mask_9;
      4'b1010 : _zz_PmpPlugin_iGuard_hits_8 = PmpPlugin_mask_10;
      4'b1011 : _zz_PmpPlugin_iGuard_hits_8 = PmpPlugin_mask_11;
      4'b1100 : _zz_PmpPlugin_iGuard_hits_8 = PmpPlugin_mask_12;
      4'b1101 : _zz_PmpPlugin_iGuard_hits_8 = PmpPlugin_mask_13;
      4'b1110 : _zz_PmpPlugin_iGuard_hits_8 = PmpPlugin_mask_14;
      default : _zz_PmpPlugin_iGuard_hits_8 = PmpPlugin_mask_15;
    endcase
  end

  always @(*) begin
    case(_zz_PmpPlugin_iGuard_hits_8_3)
      4'b0000 : _zz_PmpPlugin_iGuard_hits_8_2 = PmpPlugin_base_0;
      4'b0001 : _zz_PmpPlugin_iGuard_hits_8_2 = PmpPlugin_base_1;
      4'b0010 : _zz_PmpPlugin_iGuard_hits_8_2 = PmpPlugin_base_2;
      4'b0011 : _zz_PmpPlugin_iGuard_hits_8_2 = PmpPlugin_base_3;
      4'b0100 : _zz_PmpPlugin_iGuard_hits_8_2 = PmpPlugin_base_4;
      4'b0101 : _zz_PmpPlugin_iGuard_hits_8_2 = PmpPlugin_base_5;
      4'b0110 : _zz_PmpPlugin_iGuard_hits_8_2 = PmpPlugin_base_6;
      4'b0111 : _zz_PmpPlugin_iGuard_hits_8_2 = PmpPlugin_base_7;
      4'b1000 : _zz_PmpPlugin_iGuard_hits_8_2 = PmpPlugin_base_8;
      4'b1001 : _zz_PmpPlugin_iGuard_hits_8_2 = PmpPlugin_base_9;
      4'b1010 : _zz_PmpPlugin_iGuard_hits_8_2 = PmpPlugin_base_10;
      4'b1011 : _zz_PmpPlugin_iGuard_hits_8_2 = PmpPlugin_base_11;
      4'b1100 : _zz_PmpPlugin_iGuard_hits_8_2 = PmpPlugin_base_12;
      4'b1101 : _zz_PmpPlugin_iGuard_hits_8_2 = PmpPlugin_base_13;
      4'b1110 : _zz_PmpPlugin_iGuard_hits_8_2 = PmpPlugin_base_14;
      default : _zz_PmpPlugin_iGuard_hits_8_2 = PmpPlugin_base_15;
    endcase
  end

  always @(*) begin
    case(_zz_PmpPlugin_iGuard_hits_9_1)
      4'b0000 : _zz_PmpPlugin_iGuard_hits_9 = PmpPlugin_mask_0;
      4'b0001 : _zz_PmpPlugin_iGuard_hits_9 = PmpPlugin_mask_1;
      4'b0010 : _zz_PmpPlugin_iGuard_hits_9 = PmpPlugin_mask_2;
      4'b0011 : _zz_PmpPlugin_iGuard_hits_9 = PmpPlugin_mask_3;
      4'b0100 : _zz_PmpPlugin_iGuard_hits_9 = PmpPlugin_mask_4;
      4'b0101 : _zz_PmpPlugin_iGuard_hits_9 = PmpPlugin_mask_5;
      4'b0110 : _zz_PmpPlugin_iGuard_hits_9 = PmpPlugin_mask_6;
      4'b0111 : _zz_PmpPlugin_iGuard_hits_9 = PmpPlugin_mask_7;
      4'b1000 : _zz_PmpPlugin_iGuard_hits_9 = PmpPlugin_mask_8;
      4'b1001 : _zz_PmpPlugin_iGuard_hits_9 = PmpPlugin_mask_9;
      4'b1010 : _zz_PmpPlugin_iGuard_hits_9 = PmpPlugin_mask_10;
      4'b1011 : _zz_PmpPlugin_iGuard_hits_9 = PmpPlugin_mask_11;
      4'b1100 : _zz_PmpPlugin_iGuard_hits_9 = PmpPlugin_mask_12;
      4'b1101 : _zz_PmpPlugin_iGuard_hits_9 = PmpPlugin_mask_13;
      4'b1110 : _zz_PmpPlugin_iGuard_hits_9 = PmpPlugin_mask_14;
      default : _zz_PmpPlugin_iGuard_hits_9 = PmpPlugin_mask_15;
    endcase
  end

  always @(*) begin
    case(_zz_PmpPlugin_iGuard_hits_9_3)
      4'b0000 : _zz_PmpPlugin_iGuard_hits_9_2 = PmpPlugin_base_0;
      4'b0001 : _zz_PmpPlugin_iGuard_hits_9_2 = PmpPlugin_base_1;
      4'b0010 : _zz_PmpPlugin_iGuard_hits_9_2 = PmpPlugin_base_2;
      4'b0011 : _zz_PmpPlugin_iGuard_hits_9_2 = PmpPlugin_base_3;
      4'b0100 : _zz_PmpPlugin_iGuard_hits_9_2 = PmpPlugin_base_4;
      4'b0101 : _zz_PmpPlugin_iGuard_hits_9_2 = PmpPlugin_base_5;
      4'b0110 : _zz_PmpPlugin_iGuard_hits_9_2 = PmpPlugin_base_6;
      4'b0111 : _zz_PmpPlugin_iGuard_hits_9_2 = PmpPlugin_base_7;
      4'b1000 : _zz_PmpPlugin_iGuard_hits_9_2 = PmpPlugin_base_8;
      4'b1001 : _zz_PmpPlugin_iGuard_hits_9_2 = PmpPlugin_base_9;
      4'b1010 : _zz_PmpPlugin_iGuard_hits_9_2 = PmpPlugin_base_10;
      4'b1011 : _zz_PmpPlugin_iGuard_hits_9_2 = PmpPlugin_base_11;
      4'b1100 : _zz_PmpPlugin_iGuard_hits_9_2 = PmpPlugin_base_12;
      4'b1101 : _zz_PmpPlugin_iGuard_hits_9_2 = PmpPlugin_base_13;
      4'b1110 : _zz_PmpPlugin_iGuard_hits_9_2 = PmpPlugin_base_14;
      default : _zz_PmpPlugin_iGuard_hits_9_2 = PmpPlugin_base_15;
    endcase
  end

  always @(*) begin
    case(_zz_PmpPlugin_iGuard_hits_10_1)
      4'b0000 : _zz_PmpPlugin_iGuard_hits_10 = PmpPlugin_mask_0;
      4'b0001 : _zz_PmpPlugin_iGuard_hits_10 = PmpPlugin_mask_1;
      4'b0010 : _zz_PmpPlugin_iGuard_hits_10 = PmpPlugin_mask_2;
      4'b0011 : _zz_PmpPlugin_iGuard_hits_10 = PmpPlugin_mask_3;
      4'b0100 : _zz_PmpPlugin_iGuard_hits_10 = PmpPlugin_mask_4;
      4'b0101 : _zz_PmpPlugin_iGuard_hits_10 = PmpPlugin_mask_5;
      4'b0110 : _zz_PmpPlugin_iGuard_hits_10 = PmpPlugin_mask_6;
      4'b0111 : _zz_PmpPlugin_iGuard_hits_10 = PmpPlugin_mask_7;
      4'b1000 : _zz_PmpPlugin_iGuard_hits_10 = PmpPlugin_mask_8;
      4'b1001 : _zz_PmpPlugin_iGuard_hits_10 = PmpPlugin_mask_9;
      4'b1010 : _zz_PmpPlugin_iGuard_hits_10 = PmpPlugin_mask_10;
      4'b1011 : _zz_PmpPlugin_iGuard_hits_10 = PmpPlugin_mask_11;
      4'b1100 : _zz_PmpPlugin_iGuard_hits_10 = PmpPlugin_mask_12;
      4'b1101 : _zz_PmpPlugin_iGuard_hits_10 = PmpPlugin_mask_13;
      4'b1110 : _zz_PmpPlugin_iGuard_hits_10 = PmpPlugin_mask_14;
      default : _zz_PmpPlugin_iGuard_hits_10 = PmpPlugin_mask_15;
    endcase
  end

  always @(*) begin
    case(_zz_PmpPlugin_iGuard_hits_10_3)
      4'b0000 : _zz_PmpPlugin_iGuard_hits_10_2 = PmpPlugin_base_0;
      4'b0001 : _zz_PmpPlugin_iGuard_hits_10_2 = PmpPlugin_base_1;
      4'b0010 : _zz_PmpPlugin_iGuard_hits_10_2 = PmpPlugin_base_2;
      4'b0011 : _zz_PmpPlugin_iGuard_hits_10_2 = PmpPlugin_base_3;
      4'b0100 : _zz_PmpPlugin_iGuard_hits_10_2 = PmpPlugin_base_4;
      4'b0101 : _zz_PmpPlugin_iGuard_hits_10_2 = PmpPlugin_base_5;
      4'b0110 : _zz_PmpPlugin_iGuard_hits_10_2 = PmpPlugin_base_6;
      4'b0111 : _zz_PmpPlugin_iGuard_hits_10_2 = PmpPlugin_base_7;
      4'b1000 : _zz_PmpPlugin_iGuard_hits_10_2 = PmpPlugin_base_8;
      4'b1001 : _zz_PmpPlugin_iGuard_hits_10_2 = PmpPlugin_base_9;
      4'b1010 : _zz_PmpPlugin_iGuard_hits_10_2 = PmpPlugin_base_10;
      4'b1011 : _zz_PmpPlugin_iGuard_hits_10_2 = PmpPlugin_base_11;
      4'b1100 : _zz_PmpPlugin_iGuard_hits_10_2 = PmpPlugin_base_12;
      4'b1101 : _zz_PmpPlugin_iGuard_hits_10_2 = PmpPlugin_base_13;
      4'b1110 : _zz_PmpPlugin_iGuard_hits_10_2 = PmpPlugin_base_14;
      default : _zz_PmpPlugin_iGuard_hits_10_2 = PmpPlugin_base_15;
    endcase
  end

  always @(*) begin
    case(_zz_PmpPlugin_iGuard_hits_11_1)
      4'b0000 : _zz_PmpPlugin_iGuard_hits_11 = PmpPlugin_mask_0;
      4'b0001 : _zz_PmpPlugin_iGuard_hits_11 = PmpPlugin_mask_1;
      4'b0010 : _zz_PmpPlugin_iGuard_hits_11 = PmpPlugin_mask_2;
      4'b0011 : _zz_PmpPlugin_iGuard_hits_11 = PmpPlugin_mask_3;
      4'b0100 : _zz_PmpPlugin_iGuard_hits_11 = PmpPlugin_mask_4;
      4'b0101 : _zz_PmpPlugin_iGuard_hits_11 = PmpPlugin_mask_5;
      4'b0110 : _zz_PmpPlugin_iGuard_hits_11 = PmpPlugin_mask_6;
      4'b0111 : _zz_PmpPlugin_iGuard_hits_11 = PmpPlugin_mask_7;
      4'b1000 : _zz_PmpPlugin_iGuard_hits_11 = PmpPlugin_mask_8;
      4'b1001 : _zz_PmpPlugin_iGuard_hits_11 = PmpPlugin_mask_9;
      4'b1010 : _zz_PmpPlugin_iGuard_hits_11 = PmpPlugin_mask_10;
      4'b1011 : _zz_PmpPlugin_iGuard_hits_11 = PmpPlugin_mask_11;
      4'b1100 : _zz_PmpPlugin_iGuard_hits_11 = PmpPlugin_mask_12;
      4'b1101 : _zz_PmpPlugin_iGuard_hits_11 = PmpPlugin_mask_13;
      4'b1110 : _zz_PmpPlugin_iGuard_hits_11 = PmpPlugin_mask_14;
      default : _zz_PmpPlugin_iGuard_hits_11 = PmpPlugin_mask_15;
    endcase
  end

  always @(*) begin
    case(_zz_PmpPlugin_iGuard_hits_11_3)
      4'b0000 : _zz_PmpPlugin_iGuard_hits_11_2 = PmpPlugin_base_0;
      4'b0001 : _zz_PmpPlugin_iGuard_hits_11_2 = PmpPlugin_base_1;
      4'b0010 : _zz_PmpPlugin_iGuard_hits_11_2 = PmpPlugin_base_2;
      4'b0011 : _zz_PmpPlugin_iGuard_hits_11_2 = PmpPlugin_base_3;
      4'b0100 : _zz_PmpPlugin_iGuard_hits_11_2 = PmpPlugin_base_4;
      4'b0101 : _zz_PmpPlugin_iGuard_hits_11_2 = PmpPlugin_base_5;
      4'b0110 : _zz_PmpPlugin_iGuard_hits_11_2 = PmpPlugin_base_6;
      4'b0111 : _zz_PmpPlugin_iGuard_hits_11_2 = PmpPlugin_base_7;
      4'b1000 : _zz_PmpPlugin_iGuard_hits_11_2 = PmpPlugin_base_8;
      4'b1001 : _zz_PmpPlugin_iGuard_hits_11_2 = PmpPlugin_base_9;
      4'b1010 : _zz_PmpPlugin_iGuard_hits_11_2 = PmpPlugin_base_10;
      4'b1011 : _zz_PmpPlugin_iGuard_hits_11_2 = PmpPlugin_base_11;
      4'b1100 : _zz_PmpPlugin_iGuard_hits_11_2 = PmpPlugin_base_12;
      4'b1101 : _zz_PmpPlugin_iGuard_hits_11_2 = PmpPlugin_base_13;
      4'b1110 : _zz_PmpPlugin_iGuard_hits_11_2 = PmpPlugin_base_14;
      default : _zz_PmpPlugin_iGuard_hits_11_2 = PmpPlugin_base_15;
    endcase
  end

  always @(*) begin
    case(_zz_PmpPlugin_iGuard_hits_12_1)
      4'b0000 : _zz_PmpPlugin_iGuard_hits_12 = PmpPlugin_mask_0;
      4'b0001 : _zz_PmpPlugin_iGuard_hits_12 = PmpPlugin_mask_1;
      4'b0010 : _zz_PmpPlugin_iGuard_hits_12 = PmpPlugin_mask_2;
      4'b0011 : _zz_PmpPlugin_iGuard_hits_12 = PmpPlugin_mask_3;
      4'b0100 : _zz_PmpPlugin_iGuard_hits_12 = PmpPlugin_mask_4;
      4'b0101 : _zz_PmpPlugin_iGuard_hits_12 = PmpPlugin_mask_5;
      4'b0110 : _zz_PmpPlugin_iGuard_hits_12 = PmpPlugin_mask_6;
      4'b0111 : _zz_PmpPlugin_iGuard_hits_12 = PmpPlugin_mask_7;
      4'b1000 : _zz_PmpPlugin_iGuard_hits_12 = PmpPlugin_mask_8;
      4'b1001 : _zz_PmpPlugin_iGuard_hits_12 = PmpPlugin_mask_9;
      4'b1010 : _zz_PmpPlugin_iGuard_hits_12 = PmpPlugin_mask_10;
      4'b1011 : _zz_PmpPlugin_iGuard_hits_12 = PmpPlugin_mask_11;
      4'b1100 : _zz_PmpPlugin_iGuard_hits_12 = PmpPlugin_mask_12;
      4'b1101 : _zz_PmpPlugin_iGuard_hits_12 = PmpPlugin_mask_13;
      4'b1110 : _zz_PmpPlugin_iGuard_hits_12 = PmpPlugin_mask_14;
      default : _zz_PmpPlugin_iGuard_hits_12 = PmpPlugin_mask_15;
    endcase
  end

  always @(*) begin
    case(_zz_PmpPlugin_iGuard_hits_12_3)
      4'b0000 : _zz_PmpPlugin_iGuard_hits_12_2 = PmpPlugin_base_0;
      4'b0001 : _zz_PmpPlugin_iGuard_hits_12_2 = PmpPlugin_base_1;
      4'b0010 : _zz_PmpPlugin_iGuard_hits_12_2 = PmpPlugin_base_2;
      4'b0011 : _zz_PmpPlugin_iGuard_hits_12_2 = PmpPlugin_base_3;
      4'b0100 : _zz_PmpPlugin_iGuard_hits_12_2 = PmpPlugin_base_4;
      4'b0101 : _zz_PmpPlugin_iGuard_hits_12_2 = PmpPlugin_base_5;
      4'b0110 : _zz_PmpPlugin_iGuard_hits_12_2 = PmpPlugin_base_6;
      4'b0111 : _zz_PmpPlugin_iGuard_hits_12_2 = PmpPlugin_base_7;
      4'b1000 : _zz_PmpPlugin_iGuard_hits_12_2 = PmpPlugin_base_8;
      4'b1001 : _zz_PmpPlugin_iGuard_hits_12_2 = PmpPlugin_base_9;
      4'b1010 : _zz_PmpPlugin_iGuard_hits_12_2 = PmpPlugin_base_10;
      4'b1011 : _zz_PmpPlugin_iGuard_hits_12_2 = PmpPlugin_base_11;
      4'b1100 : _zz_PmpPlugin_iGuard_hits_12_2 = PmpPlugin_base_12;
      4'b1101 : _zz_PmpPlugin_iGuard_hits_12_2 = PmpPlugin_base_13;
      4'b1110 : _zz_PmpPlugin_iGuard_hits_12_2 = PmpPlugin_base_14;
      default : _zz_PmpPlugin_iGuard_hits_12_2 = PmpPlugin_base_15;
    endcase
  end

  always @(*) begin
    case(_zz_PmpPlugin_iGuard_hits_13_1)
      4'b0000 : _zz_PmpPlugin_iGuard_hits_13 = PmpPlugin_mask_0;
      4'b0001 : _zz_PmpPlugin_iGuard_hits_13 = PmpPlugin_mask_1;
      4'b0010 : _zz_PmpPlugin_iGuard_hits_13 = PmpPlugin_mask_2;
      4'b0011 : _zz_PmpPlugin_iGuard_hits_13 = PmpPlugin_mask_3;
      4'b0100 : _zz_PmpPlugin_iGuard_hits_13 = PmpPlugin_mask_4;
      4'b0101 : _zz_PmpPlugin_iGuard_hits_13 = PmpPlugin_mask_5;
      4'b0110 : _zz_PmpPlugin_iGuard_hits_13 = PmpPlugin_mask_6;
      4'b0111 : _zz_PmpPlugin_iGuard_hits_13 = PmpPlugin_mask_7;
      4'b1000 : _zz_PmpPlugin_iGuard_hits_13 = PmpPlugin_mask_8;
      4'b1001 : _zz_PmpPlugin_iGuard_hits_13 = PmpPlugin_mask_9;
      4'b1010 : _zz_PmpPlugin_iGuard_hits_13 = PmpPlugin_mask_10;
      4'b1011 : _zz_PmpPlugin_iGuard_hits_13 = PmpPlugin_mask_11;
      4'b1100 : _zz_PmpPlugin_iGuard_hits_13 = PmpPlugin_mask_12;
      4'b1101 : _zz_PmpPlugin_iGuard_hits_13 = PmpPlugin_mask_13;
      4'b1110 : _zz_PmpPlugin_iGuard_hits_13 = PmpPlugin_mask_14;
      default : _zz_PmpPlugin_iGuard_hits_13 = PmpPlugin_mask_15;
    endcase
  end

  always @(*) begin
    case(_zz_PmpPlugin_iGuard_hits_13_3)
      4'b0000 : _zz_PmpPlugin_iGuard_hits_13_2 = PmpPlugin_base_0;
      4'b0001 : _zz_PmpPlugin_iGuard_hits_13_2 = PmpPlugin_base_1;
      4'b0010 : _zz_PmpPlugin_iGuard_hits_13_2 = PmpPlugin_base_2;
      4'b0011 : _zz_PmpPlugin_iGuard_hits_13_2 = PmpPlugin_base_3;
      4'b0100 : _zz_PmpPlugin_iGuard_hits_13_2 = PmpPlugin_base_4;
      4'b0101 : _zz_PmpPlugin_iGuard_hits_13_2 = PmpPlugin_base_5;
      4'b0110 : _zz_PmpPlugin_iGuard_hits_13_2 = PmpPlugin_base_6;
      4'b0111 : _zz_PmpPlugin_iGuard_hits_13_2 = PmpPlugin_base_7;
      4'b1000 : _zz_PmpPlugin_iGuard_hits_13_2 = PmpPlugin_base_8;
      4'b1001 : _zz_PmpPlugin_iGuard_hits_13_2 = PmpPlugin_base_9;
      4'b1010 : _zz_PmpPlugin_iGuard_hits_13_2 = PmpPlugin_base_10;
      4'b1011 : _zz_PmpPlugin_iGuard_hits_13_2 = PmpPlugin_base_11;
      4'b1100 : _zz_PmpPlugin_iGuard_hits_13_2 = PmpPlugin_base_12;
      4'b1101 : _zz_PmpPlugin_iGuard_hits_13_2 = PmpPlugin_base_13;
      4'b1110 : _zz_PmpPlugin_iGuard_hits_13_2 = PmpPlugin_base_14;
      default : _zz_PmpPlugin_iGuard_hits_13_2 = PmpPlugin_base_15;
    endcase
  end

  always @(*) begin
    case(_zz_PmpPlugin_iGuard_hits_14_1)
      4'b0000 : _zz_PmpPlugin_iGuard_hits_14 = PmpPlugin_mask_0;
      4'b0001 : _zz_PmpPlugin_iGuard_hits_14 = PmpPlugin_mask_1;
      4'b0010 : _zz_PmpPlugin_iGuard_hits_14 = PmpPlugin_mask_2;
      4'b0011 : _zz_PmpPlugin_iGuard_hits_14 = PmpPlugin_mask_3;
      4'b0100 : _zz_PmpPlugin_iGuard_hits_14 = PmpPlugin_mask_4;
      4'b0101 : _zz_PmpPlugin_iGuard_hits_14 = PmpPlugin_mask_5;
      4'b0110 : _zz_PmpPlugin_iGuard_hits_14 = PmpPlugin_mask_6;
      4'b0111 : _zz_PmpPlugin_iGuard_hits_14 = PmpPlugin_mask_7;
      4'b1000 : _zz_PmpPlugin_iGuard_hits_14 = PmpPlugin_mask_8;
      4'b1001 : _zz_PmpPlugin_iGuard_hits_14 = PmpPlugin_mask_9;
      4'b1010 : _zz_PmpPlugin_iGuard_hits_14 = PmpPlugin_mask_10;
      4'b1011 : _zz_PmpPlugin_iGuard_hits_14 = PmpPlugin_mask_11;
      4'b1100 : _zz_PmpPlugin_iGuard_hits_14 = PmpPlugin_mask_12;
      4'b1101 : _zz_PmpPlugin_iGuard_hits_14 = PmpPlugin_mask_13;
      4'b1110 : _zz_PmpPlugin_iGuard_hits_14 = PmpPlugin_mask_14;
      default : _zz_PmpPlugin_iGuard_hits_14 = PmpPlugin_mask_15;
    endcase
  end

  always @(*) begin
    case(_zz_PmpPlugin_iGuard_hits_14_3)
      4'b0000 : _zz_PmpPlugin_iGuard_hits_14_2 = PmpPlugin_base_0;
      4'b0001 : _zz_PmpPlugin_iGuard_hits_14_2 = PmpPlugin_base_1;
      4'b0010 : _zz_PmpPlugin_iGuard_hits_14_2 = PmpPlugin_base_2;
      4'b0011 : _zz_PmpPlugin_iGuard_hits_14_2 = PmpPlugin_base_3;
      4'b0100 : _zz_PmpPlugin_iGuard_hits_14_2 = PmpPlugin_base_4;
      4'b0101 : _zz_PmpPlugin_iGuard_hits_14_2 = PmpPlugin_base_5;
      4'b0110 : _zz_PmpPlugin_iGuard_hits_14_2 = PmpPlugin_base_6;
      4'b0111 : _zz_PmpPlugin_iGuard_hits_14_2 = PmpPlugin_base_7;
      4'b1000 : _zz_PmpPlugin_iGuard_hits_14_2 = PmpPlugin_base_8;
      4'b1001 : _zz_PmpPlugin_iGuard_hits_14_2 = PmpPlugin_base_9;
      4'b1010 : _zz_PmpPlugin_iGuard_hits_14_2 = PmpPlugin_base_10;
      4'b1011 : _zz_PmpPlugin_iGuard_hits_14_2 = PmpPlugin_base_11;
      4'b1100 : _zz_PmpPlugin_iGuard_hits_14_2 = PmpPlugin_base_12;
      4'b1101 : _zz_PmpPlugin_iGuard_hits_14_2 = PmpPlugin_base_13;
      4'b1110 : _zz_PmpPlugin_iGuard_hits_14_2 = PmpPlugin_base_14;
      default : _zz_PmpPlugin_iGuard_hits_14_2 = PmpPlugin_base_15;
    endcase
  end

  always @(*) begin
    case(_zz_PmpPlugin_iGuard_hits_15_1)
      4'b0000 : _zz_PmpPlugin_iGuard_hits_15 = PmpPlugin_mask_0;
      4'b0001 : _zz_PmpPlugin_iGuard_hits_15 = PmpPlugin_mask_1;
      4'b0010 : _zz_PmpPlugin_iGuard_hits_15 = PmpPlugin_mask_2;
      4'b0011 : _zz_PmpPlugin_iGuard_hits_15 = PmpPlugin_mask_3;
      4'b0100 : _zz_PmpPlugin_iGuard_hits_15 = PmpPlugin_mask_4;
      4'b0101 : _zz_PmpPlugin_iGuard_hits_15 = PmpPlugin_mask_5;
      4'b0110 : _zz_PmpPlugin_iGuard_hits_15 = PmpPlugin_mask_6;
      4'b0111 : _zz_PmpPlugin_iGuard_hits_15 = PmpPlugin_mask_7;
      4'b1000 : _zz_PmpPlugin_iGuard_hits_15 = PmpPlugin_mask_8;
      4'b1001 : _zz_PmpPlugin_iGuard_hits_15 = PmpPlugin_mask_9;
      4'b1010 : _zz_PmpPlugin_iGuard_hits_15 = PmpPlugin_mask_10;
      4'b1011 : _zz_PmpPlugin_iGuard_hits_15 = PmpPlugin_mask_11;
      4'b1100 : _zz_PmpPlugin_iGuard_hits_15 = PmpPlugin_mask_12;
      4'b1101 : _zz_PmpPlugin_iGuard_hits_15 = PmpPlugin_mask_13;
      4'b1110 : _zz_PmpPlugin_iGuard_hits_15 = PmpPlugin_mask_14;
      default : _zz_PmpPlugin_iGuard_hits_15 = PmpPlugin_mask_15;
    endcase
  end

  always @(*) begin
    case(_zz_PmpPlugin_iGuard_hits_15_3)
      4'b0000 : _zz_PmpPlugin_iGuard_hits_15_2 = PmpPlugin_base_0;
      4'b0001 : _zz_PmpPlugin_iGuard_hits_15_2 = PmpPlugin_base_1;
      4'b0010 : _zz_PmpPlugin_iGuard_hits_15_2 = PmpPlugin_base_2;
      4'b0011 : _zz_PmpPlugin_iGuard_hits_15_2 = PmpPlugin_base_3;
      4'b0100 : _zz_PmpPlugin_iGuard_hits_15_2 = PmpPlugin_base_4;
      4'b0101 : _zz_PmpPlugin_iGuard_hits_15_2 = PmpPlugin_base_5;
      4'b0110 : _zz_PmpPlugin_iGuard_hits_15_2 = PmpPlugin_base_6;
      4'b0111 : _zz_PmpPlugin_iGuard_hits_15_2 = PmpPlugin_base_7;
      4'b1000 : _zz_PmpPlugin_iGuard_hits_15_2 = PmpPlugin_base_8;
      4'b1001 : _zz_PmpPlugin_iGuard_hits_15_2 = PmpPlugin_base_9;
      4'b1010 : _zz_PmpPlugin_iGuard_hits_15_2 = PmpPlugin_base_10;
      4'b1011 : _zz_PmpPlugin_iGuard_hits_15_2 = PmpPlugin_base_11;
      4'b1100 : _zz_PmpPlugin_iGuard_hits_15_2 = PmpPlugin_base_12;
      4'b1101 : _zz_PmpPlugin_iGuard_hits_15_2 = PmpPlugin_base_13;
      4'b1110 : _zz_PmpPlugin_iGuard_hits_15_2 = PmpPlugin_base_14;
      default : _zz_PmpPlugin_iGuard_hits_15_2 = PmpPlugin_base_15;
    endcase
  end

  always @(*) begin
    case(_zz_IBusCachedPlugin_mmuBus_rsp_allowExecute_18)
      4'b0000 : _zz_IBusCachedPlugin_mmuBus_rsp_allowExecute_17 = PmpPlugin_pmpcfg_0[2];
      4'b0001 : _zz_IBusCachedPlugin_mmuBus_rsp_allowExecute_17 = PmpPlugin_pmpcfg_1[2];
      4'b0010 : _zz_IBusCachedPlugin_mmuBus_rsp_allowExecute_17 = PmpPlugin_pmpcfg_2[2];
      4'b0011 : _zz_IBusCachedPlugin_mmuBus_rsp_allowExecute_17 = PmpPlugin_pmpcfg_3[2];
      4'b0100 : _zz_IBusCachedPlugin_mmuBus_rsp_allowExecute_17 = PmpPlugin_pmpcfg_4[2];
      4'b0101 : _zz_IBusCachedPlugin_mmuBus_rsp_allowExecute_17 = PmpPlugin_pmpcfg_5[2];
      4'b0110 : _zz_IBusCachedPlugin_mmuBus_rsp_allowExecute_17 = PmpPlugin_pmpcfg_6[2];
      4'b0111 : _zz_IBusCachedPlugin_mmuBus_rsp_allowExecute_17 = PmpPlugin_pmpcfg_7[2];
      4'b1000 : _zz_IBusCachedPlugin_mmuBus_rsp_allowExecute_17 = PmpPlugin_pmpcfg_8[2];
      4'b1001 : _zz_IBusCachedPlugin_mmuBus_rsp_allowExecute_17 = PmpPlugin_pmpcfg_9[2];
      4'b1010 : _zz_IBusCachedPlugin_mmuBus_rsp_allowExecute_17 = PmpPlugin_pmpcfg_10[2];
      4'b1011 : _zz_IBusCachedPlugin_mmuBus_rsp_allowExecute_17 = PmpPlugin_pmpcfg_11[2];
      4'b1100 : _zz_IBusCachedPlugin_mmuBus_rsp_allowExecute_17 = PmpPlugin_pmpcfg_12[2];
      4'b1101 : _zz_IBusCachedPlugin_mmuBus_rsp_allowExecute_17 = PmpPlugin_pmpcfg_13[2];
      4'b1110 : _zz_IBusCachedPlugin_mmuBus_rsp_allowExecute_17 = PmpPlugin_pmpcfg_14[2];
      default : _zz_IBusCachedPlugin_mmuBus_rsp_allowExecute_17 = PmpPlugin_pmpcfg_15[2];
    endcase
  end

  always @(*) begin
    case(_zz_when_PmpPlugin_l209_1)
      4'b0000 : _zz_when_PmpPlugin_l209 = PmpPlugin_pmpcfg_0;
      4'b0001 : _zz_when_PmpPlugin_l209 = PmpPlugin_pmpcfg_1;
      4'b0010 : _zz_when_PmpPlugin_l209 = PmpPlugin_pmpcfg_2;
      4'b0011 : _zz_when_PmpPlugin_l209 = PmpPlugin_pmpcfg_3;
      4'b0100 : _zz_when_PmpPlugin_l209 = PmpPlugin_pmpcfg_4;
      4'b0101 : _zz_when_PmpPlugin_l209 = PmpPlugin_pmpcfg_5;
      4'b0110 : _zz_when_PmpPlugin_l209 = PmpPlugin_pmpcfg_6;
      4'b0111 : _zz_when_PmpPlugin_l209 = PmpPlugin_pmpcfg_7;
      4'b1000 : _zz_when_PmpPlugin_l209 = PmpPlugin_pmpcfg_8;
      4'b1001 : _zz_when_PmpPlugin_l209 = PmpPlugin_pmpcfg_9;
      4'b1010 : _zz_when_PmpPlugin_l209 = PmpPlugin_pmpcfg_10;
      4'b1011 : _zz_when_PmpPlugin_l209 = PmpPlugin_pmpcfg_11;
      4'b1100 : _zz_when_PmpPlugin_l209 = PmpPlugin_pmpcfg_12;
      4'b1101 : _zz_when_PmpPlugin_l209 = PmpPlugin_pmpcfg_13;
      4'b1110 : _zz_when_PmpPlugin_l209 = PmpPlugin_pmpcfg_14;
      default : _zz_when_PmpPlugin_l209 = PmpPlugin_pmpcfg_15;
    endcase
  end

  always @(*) begin
    case(_zz_when_PmpPlugin_l209_1_2)
      4'b0000 : _zz_when_PmpPlugin_l209_1_1 = PmpPlugin_pmpcfg_0;
      4'b0001 : _zz_when_PmpPlugin_l209_1_1 = PmpPlugin_pmpcfg_1;
      4'b0010 : _zz_when_PmpPlugin_l209_1_1 = PmpPlugin_pmpcfg_2;
      4'b0011 : _zz_when_PmpPlugin_l209_1_1 = PmpPlugin_pmpcfg_3;
      4'b0100 : _zz_when_PmpPlugin_l209_1_1 = PmpPlugin_pmpcfg_4;
      4'b0101 : _zz_when_PmpPlugin_l209_1_1 = PmpPlugin_pmpcfg_5;
      4'b0110 : _zz_when_PmpPlugin_l209_1_1 = PmpPlugin_pmpcfg_6;
      4'b0111 : _zz_when_PmpPlugin_l209_1_1 = PmpPlugin_pmpcfg_7;
      4'b1000 : _zz_when_PmpPlugin_l209_1_1 = PmpPlugin_pmpcfg_8;
      4'b1001 : _zz_when_PmpPlugin_l209_1_1 = PmpPlugin_pmpcfg_9;
      4'b1010 : _zz_when_PmpPlugin_l209_1_1 = PmpPlugin_pmpcfg_10;
      4'b1011 : _zz_when_PmpPlugin_l209_1_1 = PmpPlugin_pmpcfg_11;
      4'b1100 : _zz_when_PmpPlugin_l209_1_1 = PmpPlugin_pmpcfg_12;
      4'b1101 : _zz_when_PmpPlugin_l209_1_1 = PmpPlugin_pmpcfg_13;
      4'b1110 : _zz_when_PmpPlugin_l209_1_1 = PmpPlugin_pmpcfg_14;
      default : _zz_when_PmpPlugin_l209_1_1 = PmpPlugin_pmpcfg_15;
    endcase
  end

  always @(*) begin
    case(_zz_when_PmpPlugin_l209_2_1)
      4'b0000 : _zz_when_PmpPlugin_l209_2 = PmpPlugin_pmpcfg_0;
      4'b0001 : _zz_when_PmpPlugin_l209_2 = PmpPlugin_pmpcfg_1;
      4'b0010 : _zz_when_PmpPlugin_l209_2 = PmpPlugin_pmpcfg_2;
      4'b0011 : _zz_when_PmpPlugin_l209_2 = PmpPlugin_pmpcfg_3;
      4'b0100 : _zz_when_PmpPlugin_l209_2 = PmpPlugin_pmpcfg_4;
      4'b0101 : _zz_when_PmpPlugin_l209_2 = PmpPlugin_pmpcfg_5;
      4'b0110 : _zz_when_PmpPlugin_l209_2 = PmpPlugin_pmpcfg_6;
      4'b0111 : _zz_when_PmpPlugin_l209_2 = PmpPlugin_pmpcfg_7;
      4'b1000 : _zz_when_PmpPlugin_l209_2 = PmpPlugin_pmpcfg_8;
      4'b1001 : _zz_when_PmpPlugin_l209_2 = PmpPlugin_pmpcfg_9;
      4'b1010 : _zz_when_PmpPlugin_l209_2 = PmpPlugin_pmpcfg_10;
      4'b1011 : _zz_when_PmpPlugin_l209_2 = PmpPlugin_pmpcfg_11;
      4'b1100 : _zz_when_PmpPlugin_l209_2 = PmpPlugin_pmpcfg_12;
      4'b1101 : _zz_when_PmpPlugin_l209_2 = PmpPlugin_pmpcfg_13;
      4'b1110 : _zz_when_PmpPlugin_l209_2 = PmpPlugin_pmpcfg_14;
      default : _zz_when_PmpPlugin_l209_2 = PmpPlugin_pmpcfg_15;
    endcase
  end

  always @(*) begin
    case(_zz_when_PmpPlugin_l209_3_1)
      4'b0000 : _zz_when_PmpPlugin_l209_3 = PmpPlugin_pmpcfg_0;
      4'b0001 : _zz_when_PmpPlugin_l209_3 = PmpPlugin_pmpcfg_1;
      4'b0010 : _zz_when_PmpPlugin_l209_3 = PmpPlugin_pmpcfg_2;
      4'b0011 : _zz_when_PmpPlugin_l209_3 = PmpPlugin_pmpcfg_3;
      4'b0100 : _zz_when_PmpPlugin_l209_3 = PmpPlugin_pmpcfg_4;
      4'b0101 : _zz_when_PmpPlugin_l209_3 = PmpPlugin_pmpcfg_5;
      4'b0110 : _zz_when_PmpPlugin_l209_3 = PmpPlugin_pmpcfg_6;
      4'b0111 : _zz_when_PmpPlugin_l209_3 = PmpPlugin_pmpcfg_7;
      4'b1000 : _zz_when_PmpPlugin_l209_3 = PmpPlugin_pmpcfg_8;
      4'b1001 : _zz_when_PmpPlugin_l209_3 = PmpPlugin_pmpcfg_9;
      4'b1010 : _zz_when_PmpPlugin_l209_3 = PmpPlugin_pmpcfg_10;
      4'b1011 : _zz_when_PmpPlugin_l209_3 = PmpPlugin_pmpcfg_11;
      4'b1100 : _zz_when_PmpPlugin_l209_3 = PmpPlugin_pmpcfg_12;
      4'b1101 : _zz_when_PmpPlugin_l209_3 = PmpPlugin_pmpcfg_13;
      4'b1110 : _zz_when_PmpPlugin_l209_3 = PmpPlugin_pmpcfg_14;
      default : _zz_when_PmpPlugin_l209_3 = PmpPlugin_pmpcfg_15;
    endcase
  end

  always @(*) begin
    case(execute_PmpPlugin_pmpNcfg_)
      4'b0000 : _zz_when_PmpPlugin_l216 = PmpPlugin_pmpcfg_0;
      4'b0001 : _zz_when_PmpPlugin_l216 = PmpPlugin_pmpcfg_1;
      4'b0010 : _zz_when_PmpPlugin_l216 = PmpPlugin_pmpcfg_2;
      4'b0011 : _zz_when_PmpPlugin_l216 = PmpPlugin_pmpcfg_3;
      4'b0100 : _zz_when_PmpPlugin_l216 = PmpPlugin_pmpcfg_4;
      4'b0101 : _zz_when_PmpPlugin_l216 = PmpPlugin_pmpcfg_5;
      4'b0110 : _zz_when_PmpPlugin_l216 = PmpPlugin_pmpcfg_6;
      4'b0111 : _zz_when_PmpPlugin_l216 = PmpPlugin_pmpcfg_7;
      4'b1000 : _zz_when_PmpPlugin_l216 = PmpPlugin_pmpcfg_8;
      4'b1001 : _zz_when_PmpPlugin_l216 = PmpPlugin_pmpcfg_9;
      4'b1010 : _zz_when_PmpPlugin_l216 = PmpPlugin_pmpcfg_10;
      4'b1011 : _zz_when_PmpPlugin_l216 = PmpPlugin_pmpcfg_11;
      4'b1100 : _zz_when_PmpPlugin_l216 = PmpPlugin_pmpcfg_12;
      4'b1101 : _zz_when_PmpPlugin_l216 = PmpPlugin_pmpcfg_13;
      4'b1110 : _zz_when_PmpPlugin_l216 = PmpPlugin_pmpcfg_14;
      default : _zz_when_PmpPlugin_l216 = PmpPlugin_pmpcfg_15;
    endcase
  end

  always @(*) begin
    case(_zz_CsrPlugin_csrMapping_readDataSignal_1)
      4'b0000 : _zz_CsrPlugin_csrMapping_readDataSignal = PmpPlugin_pmpcfg_0;
      4'b0001 : _zz_CsrPlugin_csrMapping_readDataSignal = PmpPlugin_pmpcfg_1;
      4'b0010 : _zz_CsrPlugin_csrMapping_readDataSignal = PmpPlugin_pmpcfg_2;
      4'b0011 : _zz_CsrPlugin_csrMapping_readDataSignal = PmpPlugin_pmpcfg_3;
      4'b0100 : _zz_CsrPlugin_csrMapping_readDataSignal = PmpPlugin_pmpcfg_4;
      4'b0101 : _zz_CsrPlugin_csrMapping_readDataSignal = PmpPlugin_pmpcfg_5;
      4'b0110 : _zz_CsrPlugin_csrMapping_readDataSignal = PmpPlugin_pmpcfg_6;
      4'b0111 : _zz_CsrPlugin_csrMapping_readDataSignal = PmpPlugin_pmpcfg_7;
      4'b1000 : _zz_CsrPlugin_csrMapping_readDataSignal = PmpPlugin_pmpcfg_8;
      4'b1001 : _zz_CsrPlugin_csrMapping_readDataSignal = PmpPlugin_pmpcfg_9;
      4'b1010 : _zz_CsrPlugin_csrMapping_readDataSignal = PmpPlugin_pmpcfg_10;
      4'b1011 : _zz_CsrPlugin_csrMapping_readDataSignal = PmpPlugin_pmpcfg_11;
      4'b1100 : _zz_CsrPlugin_csrMapping_readDataSignal = PmpPlugin_pmpcfg_12;
      4'b1101 : _zz_CsrPlugin_csrMapping_readDataSignal = PmpPlugin_pmpcfg_13;
      4'b1110 : _zz_CsrPlugin_csrMapping_readDataSignal = PmpPlugin_pmpcfg_14;
      default : _zz_CsrPlugin_csrMapping_readDataSignal = PmpPlugin_pmpcfg_15;
    endcase
  end

  always @(*) begin
    case(_zz_CsrPlugin_csrMapping_readDataSignal_3)
      4'b0000 : _zz_CsrPlugin_csrMapping_readDataSignal_2 = PmpPlugin_pmpcfg_0;
      4'b0001 : _zz_CsrPlugin_csrMapping_readDataSignal_2 = PmpPlugin_pmpcfg_1;
      4'b0010 : _zz_CsrPlugin_csrMapping_readDataSignal_2 = PmpPlugin_pmpcfg_2;
      4'b0011 : _zz_CsrPlugin_csrMapping_readDataSignal_2 = PmpPlugin_pmpcfg_3;
      4'b0100 : _zz_CsrPlugin_csrMapping_readDataSignal_2 = PmpPlugin_pmpcfg_4;
      4'b0101 : _zz_CsrPlugin_csrMapping_readDataSignal_2 = PmpPlugin_pmpcfg_5;
      4'b0110 : _zz_CsrPlugin_csrMapping_readDataSignal_2 = PmpPlugin_pmpcfg_6;
      4'b0111 : _zz_CsrPlugin_csrMapping_readDataSignal_2 = PmpPlugin_pmpcfg_7;
      4'b1000 : _zz_CsrPlugin_csrMapping_readDataSignal_2 = PmpPlugin_pmpcfg_8;
      4'b1001 : _zz_CsrPlugin_csrMapping_readDataSignal_2 = PmpPlugin_pmpcfg_9;
      4'b1010 : _zz_CsrPlugin_csrMapping_readDataSignal_2 = PmpPlugin_pmpcfg_10;
      4'b1011 : _zz_CsrPlugin_csrMapping_readDataSignal_2 = PmpPlugin_pmpcfg_11;
      4'b1100 : _zz_CsrPlugin_csrMapping_readDataSignal_2 = PmpPlugin_pmpcfg_12;
      4'b1101 : _zz_CsrPlugin_csrMapping_readDataSignal_2 = PmpPlugin_pmpcfg_13;
      4'b1110 : _zz_CsrPlugin_csrMapping_readDataSignal_2 = PmpPlugin_pmpcfg_14;
      default : _zz_CsrPlugin_csrMapping_readDataSignal_2 = PmpPlugin_pmpcfg_15;
    endcase
  end

  always @(*) begin
    case(_zz_CsrPlugin_csrMapping_readDataSignal_5)
      4'b0000 : _zz_CsrPlugin_csrMapping_readDataSignal_4 = PmpPlugin_pmpcfg_0;
      4'b0001 : _zz_CsrPlugin_csrMapping_readDataSignal_4 = PmpPlugin_pmpcfg_1;
      4'b0010 : _zz_CsrPlugin_csrMapping_readDataSignal_4 = PmpPlugin_pmpcfg_2;
      4'b0011 : _zz_CsrPlugin_csrMapping_readDataSignal_4 = PmpPlugin_pmpcfg_3;
      4'b0100 : _zz_CsrPlugin_csrMapping_readDataSignal_4 = PmpPlugin_pmpcfg_4;
      4'b0101 : _zz_CsrPlugin_csrMapping_readDataSignal_4 = PmpPlugin_pmpcfg_5;
      4'b0110 : _zz_CsrPlugin_csrMapping_readDataSignal_4 = PmpPlugin_pmpcfg_6;
      4'b0111 : _zz_CsrPlugin_csrMapping_readDataSignal_4 = PmpPlugin_pmpcfg_7;
      4'b1000 : _zz_CsrPlugin_csrMapping_readDataSignal_4 = PmpPlugin_pmpcfg_8;
      4'b1001 : _zz_CsrPlugin_csrMapping_readDataSignal_4 = PmpPlugin_pmpcfg_9;
      4'b1010 : _zz_CsrPlugin_csrMapping_readDataSignal_4 = PmpPlugin_pmpcfg_10;
      4'b1011 : _zz_CsrPlugin_csrMapping_readDataSignal_4 = PmpPlugin_pmpcfg_11;
      4'b1100 : _zz_CsrPlugin_csrMapping_readDataSignal_4 = PmpPlugin_pmpcfg_12;
      4'b1101 : _zz_CsrPlugin_csrMapping_readDataSignal_4 = PmpPlugin_pmpcfg_13;
      4'b1110 : _zz_CsrPlugin_csrMapping_readDataSignal_4 = PmpPlugin_pmpcfg_14;
      default : _zz_CsrPlugin_csrMapping_readDataSignal_4 = PmpPlugin_pmpcfg_15;
    endcase
  end

  always @(*) begin
    case(_zz_CsrPlugin_csrMapping_readDataSignal_7)
      4'b0000 : _zz_CsrPlugin_csrMapping_readDataSignal_6 = PmpPlugin_pmpcfg_0;
      4'b0001 : _zz_CsrPlugin_csrMapping_readDataSignal_6 = PmpPlugin_pmpcfg_1;
      4'b0010 : _zz_CsrPlugin_csrMapping_readDataSignal_6 = PmpPlugin_pmpcfg_2;
      4'b0011 : _zz_CsrPlugin_csrMapping_readDataSignal_6 = PmpPlugin_pmpcfg_3;
      4'b0100 : _zz_CsrPlugin_csrMapping_readDataSignal_6 = PmpPlugin_pmpcfg_4;
      4'b0101 : _zz_CsrPlugin_csrMapping_readDataSignal_6 = PmpPlugin_pmpcfg_5;
      4'b0110 : _zz_CsrPlugin_csrMapping_readDataSignal_6 = PmpPlugin_pmpcfg_6;
      4'b0111 : _zz_CsrPlugin_csrMapping_readDataSignal_6 = PmpPlugin_pmpcfg_7;
      4'b1000 : _zz_CsrPlugin_csrMapping_readDataSignal_6 = PmpPlugin_pmpcfg_8;
      4'b1001 : _zz_CsrPlugin_csrMapping_readDataSignal_6 = PmpPlugin_pmpcfg_9;
      4'b1010 : _zz_CsrPlugin_csrMapping_readDataSignal_6 = PmpPlugin_pmpcfg_10;
      4'b1011 : _zz_CsrPlugin_csrMapping_readDataSignal_6 = PmpPlugin_pmpcfg_11;
      4'b1100 : _zz_CsrPlugin_csrMapping_readDataSignal_6 = PmpPlugin_pmpcfg_12;
      4'b1101 : _zz_CsrPlugin_csrMapping_readDataSignal_6 = PmpPlugin_pmpcfg_13;
      4'b1110 : _zz_CsrPlugin_csrMapping_readDataSignal_6 = PmpPlugin_pmpcfg_14;
      default : _zz_CsrPlugin_csrMapping_readDataSignal_6 = PmpPlugin_pmpcfg_15;
    endcase
  end

  `ifndef SYNTHESIS
  always @(*) begin
    case(_zz_memory_to_writeBack_ENV_CTRL)
      EnvCtrlEnum_NONE : _zz_memory_to_writeBack_ENV_CTRL_string = "NONE ";
      EnvCtrlEnum_XRET : _zz_memory_to_writeBack_ENV_CTRL_string = "XRET ";
      EnvCtrlEnum_WFI : _zz_memory_to_writeBack_ENV_CTRL_string = "WFI  ";
      EnvCtrlEnum_ECALL : _zz_memory_to_writeBack_ENV_CTRL_string = "ECALL";
      default : _zz_memory_to_writeBack_ENV_CTRL_string = "?????";
    endcase
  end
  always @(*) begin
    case(_zz_memory_to_writeBack_ENV_CTRL_1)
      EnvCtrlEnum_NONE : _zz_memory_to_writeBack_ENV_CTRL_1_string = "NONE ";
      EnvCtrlEnum_XRET : _zz_memory_to_writeBack_ENV_CTRL_1_string = "XRET ";
      EnvCtrlEnum_WFI : _zz_memory_to_writeBack_ENV_CTRL_1_string = "WFI  ";
      EnvCtrlEnum_ECALL : _zz_memory_to_writeBack_ENV_CTRL_1_string = "ECALL";
      default : _zz_memory_to_writeBack_ENV_CTRL_1_string = "?????";
    endcase
  end
  always @(*) begin
    case(_zz_execute_to_memory_ENV_CTRL)
      EnvCtrlEnum_NONE : _zz_execute_to_memory_ENV_CTRL_string = "NONE ";
      EnvCtrlEnum_XRET : _zz_execute_to_memory_ENV_CTRL_string = "XRET ";
      EnvCtrlEnum_WFI : _zz_execute_to_memory_ENV_CTRL_string = "WFI  ";
      EnvCtrlEnum_ECALL : _zz_execute_to_memory_ENV_CTRL_string = "ECALL";
      default : _zz_execute_to_memory_ENV_CTRL_string = "?????";
    endcase
  end
  always @(*) begin
    case(_zz_execute_to_memory_ENV_CTRL_1)
      EnvCtrlEnum_NONE : _zz_execute_to_memory_ENV_CTRL_1_string = "NONE ";
      EnvCtrlEnum_XRET : _zz_execute_to_memory_ENV_CTRL_1_string = "XRET ";
      EnvCtrlEnum_WFI : _zz_execute_to_memory_ENV_CTRL_1_string = "WFI  ";
      EnvCtrlEnum_ECALL : _zz_execute_to_memory_ENV_CTRL_1_string = "ECALL";
      default : _zz_execute_to_memory_ENV_CTRL_1_string = "?????";
    endcase
  end
  always @(*) begin
    case(decode_ENV_CTRL)
      EnvCtrlEnum_NONE : decode_ENV_CTRL_string = "NONE ";
      EnvCtrlEnum_XRET : decode_ENV_CTRL_string = "XRET ";
      EnvCtrlEnum_WFI : decode_ENV_CTRL_string = "WFI  ";
      EnvCtrlEnum_ECALL : decode_ENV_CTRL_string = "ECALL";
      default : decode_ENV_CTRL_string = "?????";
    endcase
  end
  always @(*) begin
    case(_zz_decode_ENV_CTRL)
      EnvCtrlEnum_NONE : _zz_decode_ENV_CTRL_string = "NONE ";
      EnvCtrlEnum_XRET : _zz_decode_ENV_CTRL_string = "XRET ";
      EnvCtrlEnum_WFI : _zz_decode_ENV_CTRL_string = "WFI  ";
      EnvCtrlEnum_ECALL : _zz_decode_ENV_CTRL_string = "ECALL";
      default : _zz_decode_ENV_CTRL_string = "?????";
    endcase
  end
  always @(*) begin
    case(_zz_decode_to_execute_ENV_CTRL)
      EnvCtrlEnum_NONE : _zz_decode_to_execute_ENV_CTRL_string = "NONE ";
      EnvCtrlEnum_XRET : _zz_decode_to_execute_ENV_CTRL_string = "XRET ";
      EnvCtrlEnum_WFI : _zz_decode_to_execute_ENV_CTRL_string = "WFI  ";
      EnvCtrlEnum_ECALL : _zz_decode_to_execute_ENV_CTRL_string = "ECALL";
      default : _zz_decode_to_execute_ENV_CTRL_string = "?????";
    endcase
  end
  always @(*) begin
    case(_zz_decode_to_execute_ENV_CTRL_1)
      EnvCtrlEnum_NONE : _zz_decode_to_execute_ENV_CTRL_1_string = "NONE ";
      EnvCtrlEnum_XRET : _zz_decode_to_execute_ENV_CTRL_1_string = "XRET ";
      EnvCtrlEnum_WFI : _zz_decode_to_execute_ENV_CTRL_1_string = "WFI  ";
      EnvCtrlEnum_ECALL : _zz_decode_to_execute_ENV_CTRL_1_string = "ECALL";
      default : _zz_decode_to_execute_ENV_CTRL_1_string = "?????";
    endcase
  end
  always @(*) begin
    case(_zz_decode_to_execute_BRANCH_CTRL)
      BranchCtrlEnum_INC : _zz_decode_to_execute_BRANCH_CTRL_string = "INC ";
      BranchCtrlEnum_B : _zz_decode_to_execute_BRANCH_CTRL_string = "B   ";
      BranchCtrlEnum_JAL : _zz_decode_to_execute_BRANCH_CTRL_string = "JAL ";
      BranchCtrlEnum_JALR : _zz_decode_to_execute_BRANCH_CTRL_string = "JALR";
      default : _zz_decode_to_execute_BRANCH_CTRL_string = "????";
    endcase
  end
  always @(*) begin
    case(_zz_decode_to_execute_BRANCH_CTRL_1)
      BranchCtrlEnum_INC : _zz_decode_to_execute_BRANCH_CTRL_1_string = "INC ";
      BranchCtrlEnum_B : _zz_decode_to_execute_BRANCH_CTRL_1_string = "B   ";
      BranchCtrlEnum_JAL : _zz_decode_to_execute_BRANCH_CTRL_1_string = "JAL ";
      BranchCtrlEnum_JALR : _zz_decode_to_execute_BRANCH_CTRL_1_string = "JALR";
      default : _zz_decode_to_execute_BRANCH_CTRL_1_string = "????";
    endcase
  end
  always @(*) begin
    case(_zz_execute_to_memory_SHIFT_CTRL)
      ShiftCtrlEnum_DISABLE_1 : _zz_execute_to_memory_SHIFT_CTRL_string = "DISABLE_1";
      ShiftCtrlEnum_SLL_1 : _zz_execute_to_memory_SHIFT_CTRL_string = "SLL_1    ";
      ShiftCtrlEnum_SRL_1 : _zz_execute_to_memory_SHIFT_CTRL_string = "SRL_1    ";
      ShiftCtrlEnum_SRA_1 : _zz_execute_to_memory_SHIFT_CTRL_string = "SRA_1    ";
      default : _zz_execute_to_memory_SHIFT_CTRL_string = "?????????";
    endcase
  end
  always @(*) begin
    case(_zz_execute_to_memory_SHIFT_CTRL_1)
      ShiftCtrlEnum_DISABLE_1 : _zz_execute_to_memory_SHIFT_CTRL_1_string = "DISABLE_1";
      ShiftCtrlEnum_SLL_1 : _zz_execute_to_memory_SHIFT_CTRL_1_string = "SLL_1    ";
      ShiftCtrlEnum_SRL_1 : _zz_execute_to_memory_SHIFT_CTRL_1_string = "SRL_1    ";
      ShiftCtrlEnum_SRA_1 : _zz_execute_to_memory_SHIFT_CTRL_1_string = "SRA_1    ";
      default : _zz_execute_to_memory_SHIFT_CTRL_1_string = "?????????";
    endcase
  end
  always @(*) begin
    case(decode_SHIFT_CTRL)
      ShiftCtrlEnum_DISABLE_1 : decode_SHIFT_CTRL_string = "DISABLE_1";
      ShiftCtrlEnum_SLL_1 : decode_SHIFT_CTRL_string = "SLL_1    ";
      ShiftCtrlEnum_SRL_1 : decode_SHIFT_CTRL_string = "SRL_1    ";
      ShiftCtrlEnum_SRA_1 : decode_SHIFT_CTRL_string = "SRA_1    ";
      default : decode_SHIFT_CTRL_string = "?????????";
    endcase
  end
  always @(*) begin
    case(_zz_decode_SHIFT_CTRL)
      ShiftCtrlEnum_DISABLE_1 : _zz_decode_SHIFT_CTRL_string = "DISABLE_1";
      ShiftCtrlEnum_SLL_1 : _zz_decode_SHIFT_CTRL_string = "SLL_1    ";
      ShiftCtrlEnum_SRL_1 : _zz_decode_SHIFT_CTRL_string = "SRL_1    ";
      ShiftCtrlEnum_SRA_1 : _zz_decode_SHIFT_CTRL_string = "SRA_1    ";
      default : _zz_decode_SHIFT_CTRL_string = "?????????";
    endcase
  end
  always @(*) begin
    case(_zz_decode_to_execute_SHIFT_CTRL)
      ShiftCtrlEnum_DISABLE_1 : _zz_decode_to_execute_SHIFT_CTRL_string = "DISABLE_1";
      ShiftCtrlEnum_SLL_1 : _zz_decode_to_execute_SHIFT_CTRL_string = "SLL_1    ";
      ShiftCtrlEnum_SRL_1 : _zz_decode_to_execute_SHIFT_CTRL_string = "SRL_1    ";
      ShiftCtrlEnum_SRA_1 : _zz_decode_to_execute_SHIFT_CTRL_string = "SRA_1    ";
      default : _zz_decode_to_execute_SHIFT_CTRL_string = "?????????";
    endcase
  end
  always @(*) begin
    case(_zz_decode_to_execute_SHIFT_CTRL_1)
      ShiftCtrlEnum_DISABLE_1 : _zz_decode_to_execute_SHIFT_CTRL_1_string = "DISABLE_1";
      ShiftCtrlEnum_SLL_1 : _zz_decode_to_execute_SHIFT_CTRL_1_string = "SLL_1    ";
      ShiftCtrlEnum_SRL_1 : _zz_decode_to_execute_SHIFT_CTRL_1_string = "SRL_1    ";
      ShiftCtrlEnum_SRA_1 : _zz_decode_to_execute_SHIFT_CTRL_1_string = "SRA_1    ";
      default : _zz_decode_to_execute_SHIFT_CTRL_1_string = "?????????";
    endcase
  end
  always @(*) begin
    case(decode_ALU_BITWISE_CTRL)
      AluBitwiseCtrlEnum_XOR_1 : decode_ALU_BITWISE_CTRL_string = "XOR_1";
      AluBitwiseCtrlEnum_OR_1 : decode_ALU_BITWISE_CTRL_string = "OR_1 ";
      AluBitwiseCtrlEnum_AND_1 : decode_ALU_BITWISE_CTRL_string = "AND_1";
      default : decode_ALU_BITWISE_CTRL_string = "?????";
    endcase
  end
  always @(*) begin
    case(_zz_decode_ALU_BITWISE_CTRL)
      AluBitwiseCtrlEnum_XOR_1 : _zz_decode_ALU_BITWISE_CTRL_string = "XOR_1";
      AluBitwiseCtrlEnum_OR_1 : _zz_decode_ALU_BITWISE_CTRL_string = "OR_1 ";
      AluBitwiseCtrlEnum_AND_1 : _zz_decode_ALU_BITWISE_CTRL_string = "AND_1";
      default : _zz_decode_ALU_BITWISE_CTRL_string = "?????";
    endcase
  end
  always @(*) begin
    case(_zz_decode_to_execute_ALU_BITWISE_CTRL)
      AluBitwiseCtrlEnum_XOR_1 : _zz_decode_to_execute_ALU_BITWISE_CTRL_string = "XOR_1";
      AluBitwiseCtrlEnum_OR_1 : _zz_decode_to_execute_ALU_BITWISE_CTRL_string = "OR_1 ";
      AluBitwiseCtrlEnum_AND_1 : _zz_decode_to_execute_ALU_BITWISE_CTRL_string = "AND_1";
      default : _zz_decode_to_execute_ALU_BITWISE_CTRL_string = "?????";
    endcase
  end
  always @(*) begin
    case(_zz_decode_to_execute_ALU_BITWISE_CTRL_1)
      AluBitwiseCtrlEnum_XOR_1 : _zz_decode_to_execute_ALU_BITWISE_CTRL_1_string = "XOR_1";
      AluBitwiseCtrlEnum_OR_1 : _zz_decode_to_execute_ALU_BITWISE_CTRL_1_string = "OR_1 ";
      AluBitwiseCtrlEnum_AND_1 : _zz_decode_to_execute_ALU_BITWISE_CTRL_1_string = "AND_1";
      default : _zz_decode_to_execute_ALU_BITWISE_CTRL_1_string = "?????";
    endcase
  end
  always @(*) begin
    case(decode_SRC2_CTRL)
      Src2CtrlEnum_RS : decode_SRC2_CTRL_string = "RS ";
      Src2CtrlEnum_IMI : decode_SRC2_CTRL_string = "IMI";
      Src2CtrlEnum_IMS : decode_SRC2_CTRL_string = "IMS";
      Src2CtrlEnum_PC : decode_SRC2_CTRL_string = "PC ";
      default : decode_SRC2_CTRL_string = "???";
    endcase
  end
  always @(*) begin
    case(_zz_decode_SRC2_CTRL)
      Src2CtrlEnum_RS : _zz_decode_SRC2_CTRL_string = "RS ";
      Src2CtrlEnum_IMI : _zz_decode_SRC2_CTRL_string = "IMI";
      Src2CtrlEnum_IMS : _zz_decode_SRC2_CTRL_string = "IMS";
      Src2CtrlEnum_PC : _zz_decode_SRC2_CTRL_string = "PC ";
      default : _zz_decode_SRC2_CTRL_string = "???";
    endcase
  end
  always @(*) begin
    case(_zz_decode_to_execute_SRC2_CTRL)
      Src2CtrlEnum_RS : _zz_decode_to_execute_SRC2_CTRL_string = "RS ";
      Src2CtrlEnum_IMI : _zz_decode_to_execute_SRC2_CTRL_string = "IMI";
      Src2CtrlEnum_IMS : _zz_decode_to_execute_SRC2_CTRL_string = "IMS";
      Src2CtrlEnum_PC : _zz_decode_to_execute_SRC2_CTRL_string = "PC ";
      default : _zz_decode_to_execute_SRC2_CTRL_string = "???";
    endcase
  end
  always @(*) begin
    case(_zz_decode_to_execute_SRC2_CTRL_1)
      Src2CtrlEnum_RS : _zz_decode_to_execute_SRC2_CTRL_1_string = "RS ";
      Src2CtrlEnum_IMI : _zz_decode_to_execute_SRC2_CTRL_1_string = "IMI";
      Src2CtrlEnum_IMS : _zz_decode_to_execute_SRC2_CTRL_1_string = "IMS";
      Src2CtrlEnum_PC : _zz_decode_to_execute_SRC2_CTRL_1_string = "PC ";
      default : _zz_decode_to_execute_SRC2_CTRL_1_string = "???";
    endcase
  end
  always @(*) begin
    case(decode_ALU_CTRL)
      AluCtrlEnum_ADD_SUB : decode_ALU_CTRL_string = "ADD_SUB ";
      AluCtrlEnum_SLT_SLTU : decode_ALU_CTRL_string = "SLT_SLTU";
      AluCtrlEnum_BITWISE : decode_ALU_CTRL_string = "BITWISE ";
      default : decode_ALU_CTRL_string = "????????";
    endcase
  end
  always @(*) begin
    case(_zz_decode_ALU_CTRL)
      AluCtrlEnum_ADD_SUB : _zz_decode_ALU_CTRL_string = "ADD_SUB ";
      AluCtrlEnum_SLT_SLTU : _zz_decode_ALU_CTRL_string = "SLT_SLTU";
      AluCtrlEnum_BITWISE : _zz_decode_ALU_CTRL_string = "BITWISE ";
      default : _zz_decode_ALU_CTRL_string = "????????";
    endcase
  end
  always @(*) begin
    case(_zz_decode_to_execute_ALU_CTRL)
      AluCtrlEnum_ADD_SUB : _zz_decode_to_execute_ALU_CTRL_string = "ADD_SUB ";
      AluCtrlEnum_SLT_SLTU : _zz_decode_to_execute_ALU_CTRL_string = "SLT_SLTU";
      AluCtrlEnum_BITWISE : _zz_decode_to_execute_ALU_CTRL_string = "BITWISE ";
      default : _zz_decode_to_execute_ALU_CTRL_string = "????????";
    endcase
  end
  always @(*) begin
    case(_zz_decode_to_execute_ALU_CTRL_1)
      AluCtrlEnum_ADD_SUB : _zz_decode_to_execute_ALU_CTRL_1_string = "ADD_SUB ";
      AluCtrlEnum_SLT_SLTU : _zz_decode_to_execute_ALU_CTRL_1_string = "SLT_SLTU";
      AluCtrlEnum_BITWISE : _zz_decode_to_execute_ALU_CTRL_1_string = "BITWISE ";
      default : _zz_decode_to_execute_ALU_CTRL_1_string = "????????";
    endcase
  end
  always @(*) begin
    case(decode_SRC1_CTRL)
      Src1CtrlEnum_RS : decode_SRC1_CTRL_string = "RS          ";
      Src1CtrlEnum_IMU : decode_SRC1_CTRL_string = "IMU         ";
      Src1CtrlEnum_PC_INCREMENT : decode_SRC1_CTRL_string = "PC_INCREMENT";
      Src1CtrlEnum_URS1 : decode_SRC1_CTRL_string = "URS1        ";
      default : decode_SRC1_CTRL_string = "????????????";
    endcase
  end
  always @(*) begin
    case(_zz_decode_SRC1_CTRL)
      Src1CtrlEnum_RS : _zz_decode_SRC1_CTRL_string = "RS          ";
      Src1CtrlEnum_IMU : _zz_decode_SRC1_CTRL_string = "IMU         ";
      Src1CtrlEnum_PC_INCREMENT : _zz_decode_SRC1_CTRL_string = "PC_INCREMENT";
      Src1CtrlEnum_URS1 : _zz_decode_SRC1_CTRL_string = "URS1        ";
      default : _zz_decode_SRC1_CTRL_string = "????????????";
    endcase
  end
  always @(*) begin
    case(_zz_decode_to_execute_SRC1_CTRL)
      Src1CtrlEnum_RS : _zz_decode_to_execute_SRC1_CTRL_string = "RS          ";
      Src1CtrlEnum_IMU : _zz_decode_to_execute_SRC1_CTRL_string = "IMU         ";
      Src1CtrlEnum_PC_INCREMENT : _zz_decode_to_execute_SRC1_CTRL_string = "PC_INCREMENT";
      Src1CtrlEnum_URS1 : _zz_decode_to_execute_SRC1_CTRL_string = "URS1        ";
      default : _zz_decode_to_execute_SRC1_CTRL_string = "????????????";
    endcase
  end
  always @(*) begin
    case(_zz_decode_to_execute_SRC1_CTRL_1)
      Src1CtrlEnum_RS : _zz_decode_to_execute_SRC1_CTRL_1_string = "RS          ";
      Src1CtrlEnum_IMU : _zz_decode_to_execute_SRC1_CTRL_1_string = "IMU         ";
      Src1CtrlEnum_PC_INCREMENT : _zz_decode_to_execute_SRC1_CTRL_1_string = "PC_INCREMENT";
      Src1CtrlEnum_URS1 : _zz_decode_to_execute_SRC1_CTRL_1_string = "URS1        ";
      default : _zz_decode_to_execute_SRC1_CTRL_1_string = "????????????";
    endcase
  end
  always @(*) begin
    case(memory_ENV_CTRL)
      EnvCtrlEnum_NONE : memory_ENV_CTRL_string = "NONE ";
      EnvCtrlEnum_XRET : memory_ENV_CTRL_string = "XRET ";
      EnvCtrlEnum_WFI : memory_ENV_CTRL_string = "WFI  ";
      EnvCtrlEnum_ECALL : memory_ENV_CTRL_string = "ECALL";
      default : memory_ENV_CTRL_string = "?????";
    endcase
  end
  always @(*) begin
    case(_zz_memory_ENV_CTRL)
      EnvCtrlEnum_NONE : _zz_memory_ENV_CTRL_string = "NONE ";
      EnvCtrlEnum_XRET : _zz_memory_ENV_CTRL_string = "XRET ";
      EnvCtrlEnum_WFI : _zz_memory_ENV_CTRL_string = "WFI  ";
      EnvCtrlEnum_ECALL : _zz_memory_ENV_CTRL_string = "ECALL";
      default : _zz_memory_ENV_CTRL_string = "?????";
    endcase
  end
  always @(*) begin
    case(execute_ENV_CTRL)
      EnvCtrlEnum_NONE : execute_ENV_CTRL_string = "NONE ";
      EnvCtrlEnum_XRET : execute_ENV_CTRL_string = "XRET ";
      EnvCtrlEnum_WFI : execute_ENV_CTRL_string = "WFI  ";
      EnvCtrlEnum_ECALL : execute_ENV_CTRL_string = "ECALL";
      default : execute_ENV_CTRL_string = "?????";
    endcase
  end
  always @(*) begin
    case(_zz_execute_ENV_CTRL)
      EnvCtrlEnum_NONE : _zz_execute_ENV_CTRL_string = "NONE ";
      EnvCtrlEnum_XRET : _zz_execute_ENV_CTRL_string = "XRET ";
      EnvCtrlEnum_WFI : _zz_execute_ENV_CTRL_string = "WFI  ";
      EnvCtrlEnum_ECALL : _zz_execute_ENV_CTRL_string = "ECALL";
      default : _zz_execute_ENV_CTRL_string = "?????";
    endcase
  end
  always @(*) begin
    case(writeBack_ENV_CTRL)
      EnvCtrlEnum_NONE : writeBack_ENV_CTRL_string = "NONE ";
      EnvCtrlEnum_XRET : writeBack_ENV_CTRL_string = "XRET ";
      EnvCtrlEnum_WFI : writeBack_ENV_CTRL_string = "WFI  ";
      EnvCtrlEnum_ECALL : writeBack_ENV_CTRL_string = "ECALL";
      default : writeBack_ENV_CTRL_string = "?????";
    endcase
  end
  always @(*) begin
    case(_zz_writeBack_ENV_CTRL)
      EnvCtrlEnum_NONE : _zz_writeBack_ENV_CTRL_string = "NONE ";
      EnvCtrlEnum_XRET : _zz_writeBack_ENV_CTRL_string = "XRET ";
      EnvCtrlEnum_WFI : _zz_writeBack_ENV_CTRL_string = "WFI  ";
      EnvCtrlEnum_ECALL : _zz_writeBack_ENV_CTRL_string = "ECALL";
      default : _zz_writeBack_ENV_CTRL_string = "?????";
    endcase
  end
  always @(*) begin
    case(execute_BRANCH_CTRL)
      BranchCtrlEnum_INC : execute_BRANCH_CTRL_string = "INC ";
      BranchCtrlEnum_B : execute_BRANCH_CTRL_string = "B   ";
      BranchCtrlEnum_JAL : execute_BRANCH_CTRL_string = "JAL ";
      BranchCtrlEnum_JALR : execute_BRANCH_CTRL_string = "JALR";
      default : execute_BRANCH_CTRL_string = "????";
    endcase
  end
  always @(*) begin
    case(_zz_execute_BRANCH_CTRL)
      BranchCtrlEnum_INC : _zz_execute_BRANCH_CTRL_string = "INC ";
      BranchCtrlEnum_B : _zz_execute_BRANCH_CTRL_string = "B   ";
      BranchCtrlEnum_JAL : _zz_execute_BRANCH_CTRL_string = "JAL ";
      BranchCtrlEnum_JALR : _zz_execute_BRANCH_CTRL_string = "JALR";
      default : _zz_execute_BRANCH_CTRL_string = "????";
    endcase
  end
  always @(*) begin
    case(memory_SHIFT_CTRL)
      ShiftCtrlEnum_DISABLE_1 : memory_SHIFT_CTRL_string = "DISABLE_1";
      ShiftCtrlEnum_SLL_1 : memory_SHIFT_CTRL_string = "SLL_1    ";
      ShiftCtrlEnum_SRL_1 : memory_SHIFT_CTRL_string = "SRL_1    ";
      ShiftCtrlEnum_SRA_1 : memory_SHIFT_CTRL_string = "SRA_1    ";
      default : memory_SHIFT_CTRL_string = "?????????";
    endcase
  end
  always @(*) begin
    case(_zz_memory_SHIFT_CTRL)
      ShiftCtrlEnum_DISABLE_1 : _zz_memory_SHIFT_CTRL_string = "DISABLE_1";
      ShiftCtrlEnum_SLL_1 : _zz_memory_SHIFT_CTRL_string = "SLL_1    ";
      ShiftCtrlEnum_SRL_1 : _zz_memory_SHIFT_CTRL_string = "SRL_1    ";
      ShiftCtrlEnum_SRA_1 : _zz_memory_SHIFT_CTRL_string = "SRA_1    ";
      default : _zz_memory_SHIFT_CTRL_string = "?????????";
    endcase
  end
  always @(*) begin
    case(execute_SHIFT_CTRL)
      ShiftCtrlEnum_DISABLE_1 : execute_SHIFT_CTRL_string = "DISABLE_1";
      ShiftCtrlEnum_SLL_1 : execute_SHIFT_CTRL_string = "SLL_1    ";
      ShiftCtrlEnum_SRL_1 : execute_SHIFT_CTRL_string = "SRL_1    ";
      ShiftCtrlEnum_SRA_1 : execute_SHIFT_CTRL_string = "SRA_1    ";
      default : execute_SHIFT_CTRL_string = "?????????";
    endcase
  end
  always @(*) begin
    case(_zz_execute_SHIFT_CTRL)
      ShiftCtrlEnum_DISABLE_1 : _zz_execute_SHIFT_CTRL_string = "DISABLE_1";
      ShiftCtrlEnum_SLL_1 : _zz_execute_SHIFT_CTRL_string = "SLL_1    ";
      ShiftCtrlEnum_SRL_1 : _zz_execute_SHIFT_CTRL_string = "SRL_1    ";
      ShiftCtrlEnum_SRA_1 : _zz_execute_SHIFT_CTRL_string = "SRA_1    ";
      default : _zz_execute_SHIFT_CTRL_string = "?????????";
    endcase
  end
  always @(*) begin
    case(execute_SRC2_CTRL)
      Src2CtrlEnum_RS : execute_SRC2_CTRL_string = "RS ";
      Src2CtrlEnum_IMI : execute_SRC2_CTRL_string = "IMI";
      Src2CtrlEnum_IMS : execute_SRC2_CTRL_string = "IMS";
      Src2CtrlEnum_PC : execute_SRC2_CTRL_string = "PC ";
      default : execute_SRC2_CTRL_string = "???";
    endcase
  end
  always @(*) begin
    case(_zz_execute_SRC2_CTRL)
      Src2CtrlEnum_RS : _zz_execute_SRC2_CTRL_string = "RS ";
      Src2CtrlEnum_IMI : _zz_execute_SRC2_CTRL_string = "IMI";
      Src2CtrlEnum_IMS : _zz_execute_SRC2_CTRL_string = "IMS";
      Src2CtrlEnum_PC : _zz_execute_SRC2_CTRL_string = "PC ";
      default : _zz_execute_SRC2_CTRL_string = "???";
    endcase
  end
  always @(*) begin
    case(execute_SRC1_CTRL)
      Src1CtrlEnum_RS : execute_SRC1_CTRL_string = "RS          ";
      Src1CtrlEnum_IMU : execute_SRC1_CTRL_string = "IMU         ";
      Src1CtrlEnum_PC_INCREMENT : execute_SRC1_CTRL_string = "PC_INCREMENT";
      Src1CtrlEnum_URS1 : execute_SRC1_CTRL_string = "URS1        ";
      default : execute_SRC1_CTRL_string = "????????????";
    endcase
  end
  always @(*) begin
    case(_zz_execute_SRC1_CTRL)
      Src1CtrlEnum_RS : _zz_execute_SRC1_CTRL_string = "RS          ";
      Src1CtrlEnum_IMU : _zz_execute_SRC1_CTRL_string = "IMU         ";
      Src1CtrlEnum_PC_INCREMENT : _zz_execute_SRC1_CTRL_string = "PC_INCREMENT";
      Src1CtrlEnum_URS1 : _zz_execute_SRC1_CTRL_string = "URS1        ";
      default : _zz_execute_SRC1_CTRL_string = "????????????";
    endcase
  end
  always @(*) begin
    case(execute_ALU_CTRL)
      AluCtrlEnum_ADD_SUB : execute_ALU_CTRL_string = "ADD_SUB ";
      AluCtrlEnum_SLT_SLTU : execute_ALU_CTRL_string = "SLT_SLTU";
      AluCtrlEnum_BITWISE : execute_ALU_CTRL_string = "BITWISE ";
      default : execute_ALU_CTRL_string = "????????";
    endcase
  end
  always @(*) begin
    case(_zz_execute_ALU_CTRL)
      AluCtrlEnum_ADD_SUB : _zz_execute_ALU_CTRL_string = "ADD_SUB ";
      AluCtrlEnum_SLT_SLTU : _zz_execute_ALU_CTRL_string = "SLT_SLTU";
      AluCtrlEnum_BITWISE : _zz_execute_ALU_CTRL_string = "BITWISE ";
      default : _zz_execute_ALU_CTRL_string = "????????";
    endcase
  end
  always @(*) begin
    case(execute_ALU_BITWISE_CTRL)
      AluBitwiseCtrlEnum_XOR_1 : execute_ALU_BITWISE_CTRL_string = "XOR_1";
      AluBitwiseCtrlEnum_OR_1 : execute_ALU_BITWISE_CTRL_string = "OR_1 ";
      AluBitwiseCtrlEnum_AND_1 : execute_ALU_BITWISE_CTRL_string = "AND_1";
      default : execute_ALU_BITWISE_CTRL_string = "?????";
    endcase
  end
  always @(*) begin
    case(_zz_execute_ALU_BITWISE_CTRL)
      AluBitwiseCtrlEnum_XOR_1 : _zz_execute_ALU_BITWISE_CTRL_string = "XOR_1";
      AluBitwiseCtrlEnum_OR_1 : _zz_execute_ALU_BITWISE_CTRL_string = "OR_1 ";
      AluBitwiseCtrlEnum_AND_1 : _zz_execute_ALU_BITWISE_CTRL_string = "AND_1";
      default : _zz_execute_ALU_BITWISE_CTRL_string = "?????";
    endcase
  end
  always @(*) begin
    case(_zz_decode_ENV_CTRL_1)
      EnvCtrlEnum_NONE : _zz_decode_ENV_CTRL_1_string = "NONE ";
      EnvCtrlEnum_XRET : _zz_decode_ENV_CTRL_1_string = "XRET ";
      EnvCtrlEnum_WFI : _zz_decode_ENV_CTRL_1_string = "WFI  ";
      EnvCtrlEnum_ECALL : _zz_decode_ENV_CTRL_1_string = "ECALL";
      default : _zz_decode_ENV_CTRL_1_string = "?????";
    endcase
  end
  always @(*) begin
    case(_zz_decode_BRANCH_CTRL)
      BranchCtrlEnum_INC : _zz_decode_BRANCH_CTRL_string = "INC ";
      BranchCtrlEnum_B : _zz_decode_BRANCH_CTRL_string = "B   ";
      BranchCtrlEnum_JAL : _zz_decode_BRANCH_CTRL_string = "JAL ";
      BranchCtrlEnum_JALR : _zz_decode_BRANCH_CTRL_string = "JALR";
      default : _zz_decode_BRANCH_CTRL_string = "????";
    endcase
  end
  always @(*) begin
    case(_zz_decode_SHIFT_CTRL_1)
      ShiftCtrlEnum_DISABLE_1 : _zz_decode_SHIFT_CTRL_1_string = "DISABLE_1";
      ShiftCtrlEnum_SLL_1 : _zz_decode_SHIFT_CTRL_1_string = "SLL_1    ";
      ShiftCtrlEnum_SRL_1 : _zz_decode_SHIFT_CTRL_1_string = "SRL_1    ";
      ShiftCtrlEnum_SRA_1 : _zz_decode_SHIFT_CTRL_1_string = "SRA_1    ";
      default : _zz_decode_SHIFT_CTRL_1_string = "?????????";
    endcase
  end
  always @(*) begin
    case(_zz_decode_ALU_BITWISE_CTRL_1)
      AluBitwiseCtrlEnum_XOR_1 : _zz_decode_ALU_BITWISE_CTRL_1_string = "XOR_1";
      AluBitwiseCtrlEnum_OR_1 : _zz_decode_ALU_BITWISE_CTRL_1_string = "OR_1 ";
      AluBitwiseCtrlEnum_AND_1 : _zz_decode_ALU_BITWISE_CTRL_1_string = "AND_1";
      default : _zz_decode_ALU_BITWISE_CTRL_1_string = "?????";
    endcase
  end
  always @(*) begin
    case(_zz_decode_SRC2_CTRL_1)
      Src2CtrlEnum_RS : _zz_decode_SRC2_CTRL_1_string = "RS ";
      Src2CtrlEnum_IMI : _zz_decode_SRC2_CTRL_1_string = "IMI";
      Src2CtrlEnum_IMS : _zz_decode_SRC2_CTRL_1_string = "IMS";
      Src2CtrlEnum_PC : _zz_decode_SRC2_CTRL_1_string = "PC ";
      default : _zz_decode_SRC2_CTRL_1_string = "???";
    endcase
  end
  always @(*) begin
    case(_zz_decode_ALU_CTRL_1)
      AluCtrlEnum_ADD_SUB : _zz_decode_ALU_CTRL_1_string = "ADD_SUB ";
      AluCtrlEnum_SLT_SLTU : _zz_decode_ALU_CTRL_1_string = "SLT_SLTU";
      AluCtrlEnum_BITWISE : _zz_decode_ALU_CTRL_1_string = "BITWISE ";
      default : _zz_decode_ALU_CTRL_1_string = "????????";
    endcase
  end
  always @(*) begin
    case(_zz_decode_SRC1_CTRL_1)
      Src1CtrlEnum_RS : _zz_decode_SRC1_CTRL_1_string = "RS          ";
      Src1CtrlEnum_IMU : _zz_decode_SRC1_CTRL_1_string = "IMU         ";
      Src1CtrlEnum_PC_INCREMENT : _zz_decode_SRC1_CTRL_1_string = "PC_INCREMENT";
      Src1CtrlEnum_URS1 : _zz_decode_SRC1_CTRL_1_string = "URS1        ";
      default : _zz_decode_SRC1_CTRL_1_string = "????????????";
    endcase
  end
  always @(*) begin
    case(decode_BRANCH_CTRL)
      BranchCtrlEnum_INC : decode_BRANCH_CTRL_string = "INC ";
      BranchCtrlEnum_B : decode_BRANCH_CTRL_string = "B   ";
      BranchCtrlEnum_JAL : decode_BRANCH_CTRL_string = "JAL ";
      BranchCtrlEnum_JALR : decode_BRANCH_CTRL_string = "JALR";
      default : decode_BRANCH_CTRL_string = "????";
    endcase
  end
  always @(*) begin
    case(_zz_decode_BRANCH_CTRL_1)
      BranchCtrlEnum_INC : _zz_decode_BRANCH_CTRL_1_string = "INC ";
      BranchCtrlEnum_B : _zz_decode_BRANCH_CTRL_1_string = "B   ";
      BranchCtrlEnum_JAL : _zz_decode_BRANCH_CTRL_1_string = "JAL ";
      BranchCtrlEnum_JALR : _zz_decode_BRANCH_CTRL_1_string = "JALR";
      default : _zz_decode_BRANCH_CTRL_1_string = "????";
    endcase
  end
  always @(*) begin
    case(_zz_decode_SRC1_CTRL_2)
      Src1CtrlEnum_RS : _zz_decode_SRC1_CTRL_2_string = "RS          ";
      Src1CtrlEnum_IMU : _zz_decode_SRC1_CTRL_2_string = "IMU         ";
      Src1CtrlEnum_PC_INCREMENT : _zz_decode_SRC1_CTRL_2_string = "PC_INCREMENT";
      Src1CtrlEnum_URS1 : _zz_decode_SRC1_CTRL_2_string = "URS1        ";
      default : _zz_decode_SRC1_CTRL_2_string = "????????????";
    endcase
  end
  always @(*) begin
    case(_zz_decode_ALU_CTRL_2)
      AluCtrlEnum_ADD_SUB : _zz_decode_ALU_CTRL_2_string = "ADD_SUB ";
      AluCtrlEnum_SLT_SLTU : _zz_decode_ALU_CTRL_2_string = "SLT_SLTU";
      AluCtrlEnum_BITWISE : _zz_decode_ALU_CTRL_2_string = "BITWISE ";
      default : _zz_decode_ALU_CTRL_2_string = "????????";
    endcase
  end
  always @(*) begin
    case(_zz_decode_SRC2_CTRL_2)
      Src2CtrlEnum_RS : _zz_decode_SRC2_CTRL_2_string = "RS ";
      Src2CtrlEnum_IMI : _zz_decode_SRC2_CTRL_2_string = "IMI";
      Src2CtrlEnum_IMS : _zz_decode_SRC2_CTRL_2_string = "IMS";
      Src2CtrlEnum_PC : _zz_decode_SRC2_CTRL_2_string = "PC ";
      default : _zz_decode_SRC2_CTRL_2_string = "???";
    endcase
  end
  always @(*) begin
    case(_zz_decode_ALU_BITWISE_CTRL_2)
      AluBitwiseCtrlEnum_XOR_1 : _zz_decode_ALU_BITWISE_CTRL_2_string = "XOR_1";
      AluBitwiseCtrlEnum_OR_1 : _zz_decode_ALU_BITWISE_CTRL_2_string = "OR_1 ";
      AluBitwiseCtrlEnum_AND_1 : _zz_decode_ALU_BITWISE_CTRL_2_string = "AND_1";
      default : _zz_decode_ALU_BITWISE_CTRL_2_string = "?????";
    endcase
  end
  always @(*) begin
    case(_zz_decode_SHIFT_CTRL_2)
      ShiftCtrlEnum_DISABLE_1 : _zz_decode_SHIFT_CTRL_2_string = "DISABLE_1";
      ShiftCtrlEnum_SLL_1 : _zz_decode_SHIFT_CTRL_2_string = "SLL_1    ";
      ShiftCtrlEnum_SRL_1 : _zz_decode_SHIFT_CTRL_2_string = "SRL_1    ";
      ShiftCtrlEnum_SRA_1 : _zz_decode_SHIFT_CTRL_2_string = "SRA_1    ";
      default : _zz_decode_SHIFT_CTRL_2_string = "?????????";
    endcase
  end
  always @(*) begin
    case(_zz_decode_BRANCH_CTRL_2)
      BranchCtrlEnum_INC : _zz_decode_BRANCH_CTRL_2_string = "INC ";
      BranchCtrlEnum_B : _zz_decode_BRANCH_CTRL_2_string = "B   ";
      BranchCtrlEnum_JAL : _zz_decode_BRANCH_CTRL_2_string = "JAL ";
      BranchCtrlEnum_JALR : _zz_decode_BRANCH_CTRL_2_string = "JALR";
      default : _zz_decode_BRANCH_CTRL_2_string = "????";
    endcase
  end
  always @(*) begin
    case(_zz_decode_ENV_CTRL_2)
      EnvCtrlEnum_NONE : _zz_decode_ENV_CTRL_2_string = "NONE ";
      EnvCtrlEnum_XRET : _zz_decode_ENV_CTRL_2_string = "XRET ";
      EnvCtrlEnum_WFI : _zz_decode_ENV_CTRL_2_string = "WFI  ";
      EnvCtrlEnum_ECALL : _zz_decode_ENV_CTRL_2_string = "ECALL";
      default : _zz_decode_ENV_CTRL_2_string = "?????";
    endcase
  end
  always @(*) begin
    case(decode_to_execute_SRC1_CTRL)
      Src1CtrlEnum_RS : decode_to_execute_SRC1_CTRL_string = "RS          ";
      Src1CtrlEnum_IMU : decode_to_execute_SRC1_CTRL_string = "IMU         ";
      Src1CtrlEnum_PC_INCREMENT : decode_to_execute_SRC1_CTRL_string = "PC_INCREMENT";
      Src1CtrlEnum_URS1 : decode_to_execute_SRC1_CTRL_string = "URS1        ";
      default : decode_to_execute_SRC1_CTRL_string = "????????????";
    endcase
  end
  always @(*) begin
    case(decode_to_execute_ALU_CTRL)
      AluCtrlEnum_ADD_SUB : decode_to_execute_ALU_CTRL_string = "ADD_SUB ";
      AluCtrlEnum_SLT_SLTU : decode_to_execute_ALU_CTRL_string = "SLT_SLTU";
      AluCtrlEnum_BITWISE : decode_to_execute_ALU_CTRL_string = "BITWISE ";
      default : decode_to_execute_ALU_CTRL_string = "????????";
    endcase
  end
  always @(*) begin
    case(decode_to_execute_SRC2_CTRL)
      Src2CtrlEnum_RS : decode_to_execute_SRC2_CTRL_string = "RS ";
      Src2CtrlEnum_IMI : decode_to_execute_SRC2_CTRL_string = "IMI";
      Src2CtrlEnum_IMS : decode_to_execute_SRC2_CTRL_string = "IMS";
      Src2CtrlEnum_PC : decode_to_execute_SRC2_CTRL_string = "PC ";
      default : decode_to_execute_SRC2_CTRL_string = "???";
    endcase
  end
  always @(*) begin
    case(decode_to_execute_ALU_BITWISE_CTRL)
      AluBitwiseCtrlEnum_XOR_1 : decode_to_execute_ALU_BITWISE_CTRL_string = "XOR_1";
      AluBitwiseCtrlEnum_OR_1 : decode_to_execute_ALU_BITWISE_CTRL_string = "OR_1 ";
      AluBitwiseCtrlEnum_AND_1 : decode_to_execute_ALU_BITWISE_CTRL_string = "AND_1";
      default : decode_to_execute_ALU_BITWISE_CTRL_string = "?????";
    endcase
  end
  always @(*) begin
    case(decode_to_execute_SHIFT_CTRL)
      ShiftCtrlEnum_DISABLE_1 : decode_to_execute_SHIFT_CTRL_string = "DISABLE_1";
      ShiftCtrlEnum_SLL_1 : decode_to_execute_SHIFT_CTRL_string = "SLL_1    ";
      ShiftCtrlEnum_SRL_1 : decode_to_execute_SHIFT_CTRL_string = "SRL_1    ";
      ShiftCtrlEnum_SRA_1 : decode_to_execute_SHIFT_CTRL_string = "SRA_1    ";
      default : decode_to_execute_SHIFT_CTRL_string = "?????????";
    endcase
  end
  always @(*) begin
    case(execute_to_memory_SHIFT_CTRL)
      ShiftCtrlEnum_DISABLE_1 : execute_to_memory_SHIFT_CTRL_string = "DISABLE_1";
      ShiftCtrlEnum_SLL_1 : execute_to_memory_SHIFT_CTRL_string = "SLL_1    ";
      ShiftCtrlEnum_SRL_1 : execute_to_memory_SHIFT_CTRL_string = "SRL_1    ";
      ShiftCtrlEnum_SRA_1 : execute_to_memory_SHIFT_CTRL_string = "SRA_1    ";
      default : execute_to_memory_SHIFT_CTRL_string = "?????????";
    endcase
  end
  always @(*) begin
    case(decode_to_execute_BRANCH_CTRL)
      BranchCtrlEnum_INC : decode_to_execute_BRANCH_CTRL_string = "INC ";
      BranchCtrlEnum_B : decode_to_execute_BRANCH_CTRL_string = "B   ";
      BranchCtrlEnum_JAL : decode_to_execute_BRANCH_CTRL_string = "JAL ";
      BranchCtrlEnum_JALR : decode_to_execute_BRANCH_CTRL_string = "JALR";
      default : decode_to_execute_BRANCH_CTRL_string = "????";
    endcase
  end
  always @(*) begin
    case(decode_to_execute_ENV_CTRL)
      EnvCtrlEnum_NONE : decode_to_execute_ENV_CTRL_string = "NONE ";
      EnvCtrlEnum_XRET : decode_to_execute_ENV_CTRL_string = "XRET ";
      EnvCtrlEnum_WFI : decode_to_execute_ENV_CTRL_string = "WFI  ";
      EnvCtrlEnum_ECALL : decode_to_execute_ENV_CTRL_string = "ECALL";
      default : decode_to_execute_ENV_CTRL_string = "?????";
    endcase
  end
  always @(*) begin
    case(execute_to_memory_ENV_CTRL)
      EnvCtrlEnum_NONE : execute_to_memory_ENV_CTRL_string = "NONE ";
      EnvCtrlEnum_XRET : execute_to_memory_ENV_CTRL_string = "XRET ";
      EnvCtrlEnum_WFI : execute_to_memory_ENV_CTRL_string = "WFI  ";
      EnvCtrlEnum_ECALL : execute_to_memory_ENV_CTRL_string = "ECALL";
      default : execute_to_memory_ENV_CTRL_string = "?????";
    endcase
  end
  always @(*) begin
    case(memory_to_writeBack_ENV_CTRL)
      EnvCtrlEnum_NONE : memory_to_writeBack_ENV_CTRL_string = "NONE ";
      EnvCtrlEnum_XRET : memory_to_writeBack_ENV_CTRL_string = "XRET ";
      EnvCtrlEnum_WFI : memory_to_writeBack_ENV_CTRL_string = "WFI  ";
      EnvCtrlEnum_ECALL : memory_to_writeBack_ENV_CTRL_string = "ECALL";
      default : memory_to_writeBack_ENV_CTRL_string = "?????";
    endcase
  end
  always @(*) begin
    case(execute_PmpPlugin_fsm_stateReg)
      execute_PmpPlugin_fsm_enumDef_BOOT : execute_PmpPlugin_fsm_stateReg_string = "BOOT      ";
      execute_PmpPlugin_fsm_enumDef_stateIdle : execute_PmpPlugin_fsm_stateReg_string = "stateIdle ";
      execute_PmpPlugin_fsm_enumDef_stateWrite : execute_PmpPlugin_fsm_stateReg_string = "stateWrite";
      execute_PmpPlugin_fsm_enumDef_stateCfg : execute_PmpPlugin_fsm_stateReg_string = "stateCfg  ";
      execute_PmpPlugin_fsm_enumDef_stateAddr : execute_PmpPlugin_fsm_stateReg_string = "stateAddr ";
      default : execute_PmpPlugin_fsm_stateReg_string = "??????????";
    endcase
  end
  always @(*) begin
    case(execute_PmpPlugin_fsm_stateNext)
      execute_PmpPlugin_fsm_enumDef_BOOT : execute_PmpPlugin_fsm_stateNext_string = "BOOT      ";
      execute_PmpPlugin_fsm_enumDef_stateIdle : execute_PmpPlugin_fsm_stateNext_string = "stateIdle ";
      execute_PmpPlugin_fsm_enumDef_stateWrite : execute_PmpPlugin_fsm_stateNext_string = "stateWrite";
      execute_PmpPlugin_fsm_enumDef_stateCfg : execute_PmpPlugin_fsm_stateNext_string = "stateCfg  ";
      execute_PmpPlugin_fsm_enumDef_stateAddr : execute_PmpPlugin_fsm_stateNext_string = "stateAddr ";
      default : execute_PmpPlugin_fsm_stateNext_string = "??????????";
    endcase
  end
  `endif

  always @(*) begin
    _zz_1 = 1'b0;
    case(execute_PmpPlugin_fsm_stateReg)
      execute_PmpPlugin_fsm_enumDef_stateIdle : begin
      end
      execute_PmpPlugin_fsm_enumDef_stateWrite : begin
        if(execute_PmpPlugin_pmpaddrCsr_) begin
          if(when_PmpPlugin_l216) begin
            _zz_1 = 1'b1;
          end
        end
      end
      execute_PmpPlugin_fsm_enumDef_stateCfg : begin
      end
      execute_PmpPlugin_fsm_enumDef_stateAddr : begin
      end
      default : begin
      end
    endcase
  end

  assign memory_MUL_LOW = ($signed(_zz_memory_MUL_LOW) + $signed(_zz_memory_MUL_LOW_7));
  assign memory_MUL_HH = execute_to_memory_MUL_HH;
  assign execute_MUL_HH = ($signed(execute_MulPlugin_aHigh) * $signed(execute_MulPlugin_bHigh));
  assign execute_MUL_HL = ($signed(execute_MulPlugin_aHigh) * $signed(execute_MulPlugin_bSLow));
  assign execute_MUL_LH = ($signed(execute_MulPlugin_aSLow) * $signed(execute_MulPlugin_bHigh));
  assign execute_MUL_LL = (execute_MulPlugin_aULow * execute_MulPlugin_bULow);
  assign execute_BRANCH_CALC = {execute_BranchPlugin_branchAdder[31 : 1],1'b0};
  assign execute_BRANCH_DO = ((execute_PREDICTION_HAD_BRANCHED2 != execute_BRANCH_COND_RESULT) || execute_BranchPlugin_missAlignedTarget);
  assign execute_SHIFT_RIGHT = _zz_execute_SHIFT_RIGHT;
  assign execute_REGFILE_WRITE_DATA = _zz_execute_REGFILE_WRITE_DATA;
  assign memory_MEMORY_STORE_DATA_RF = execute_to_memory_MEMORY_STORE_DATA_RF;
  assign execute_MEMORY_STORE_DATA_RF = _zz_execute_MEMORY_STORE_DATA_RF;
  assign decode_CSR_READ_OPCODE = (decode_INSTRUCTION[13 : 7] != 7'h20);
  assign decode_CSR_WRITE_OPCODE = (! (((decode_INSTRUCTION[14 : 13] == 2'b01) && (decode_INSTRUCTION[19 : 15] == 5'h0)) || ((decode_INSTRUCTION[14 : 13] == 2'b11) && (decode_INSTRUCTION[19 : 15] == 5'h0))));
  assign decode_PREDICTION_HAD_BRANCHED2 = IBusCachedPlugin_decodePrediction_cmd_hadBranch;
  assign decode_SRC2_FORCE_ZERO = (decode_SRC_ADD_ZERO && (! decode_SRC_USE_SUB_LESS));
  assign decode_IS_RS2_SIGNED = _zz_decode_IS_RS2_SIGNED[31];
  assign decode_IS_RS1_SIGNED = _zz_decode_IS_RS2_SIGNED[30];
  assign decode_IS_DIV = _zz_decode_IS_RS2_SIGNED[29];
  assign memory_IS_MUL = execute_to_memory_IS_MUL;
  assign execute_IS_MUL = decode_to_execute_IS_MUL;
  assign decode_IS_MUL = _zz_decode_IS_RS2_SIGNED[28];
  assign _zz_memory_to_writeBack_ENV_CTRL = _zz_memory_to_writeBack_ENV_CTRL_1;
  assign _zz_execute_to_memory_ENV_CTRL = _zz_execute_to_memory_ENV_CTRL_1;
  assign decode_ENV_CTRL = _zz_decode_ENV_CTRL;
  assign _zz_decode_to_execute_ENV_CTRL = _zz_decode_to_execute_ENV_CTRL_1;
  assign decode_IS_CSR = _zz_decode_IS_RS2_SIGNED[25];
  assign _zz_decode_to_execute_BRANCH_CTRL = _zz_decode_to_execute_BRANCH_CTRL_1;
  assign _zz_execute_to_memory_SHIFT_CTRL = _zz_execute_to_memory_SHIFT_CTRL_1;
  assign decode_SHIFT_CTRL = _zz_decode_SHIFT_CTRL;
  assign _zz_decode_to_execute_SHIFT_CTRL = _zz_decode_to_execute_SHIFT_CTRL_1;
  assign decode_ALU_BITWISE_CTRL = _zz_decode_ALU_BITWISE_CTRL;
  assign _zz_decode_to_execute_ALU_BITWISE_CTRL = _zz_decode_to_execute_ALU_BITWISE_CTRL_1;
  assign decode_SRC_LESS_UNSIGNED = _zz_decode_IS_RS2_SIGNED[17];
  assign decode_MEMORY_MANAGMENT = _zz_decode_IS_RS2_SIGNED[16];
  assign memory_MEMORY_WR = execute_to_memory_MEMORY_WR;
  assign decode_MEMORY_WR = _zz_decode_IS_RS2_SIGNED[13];
  assign execute_BYPASSABLE_MEMORY_STAGE = decode_to_execute_BYPASSABLE_MEMORY_STAGE;
  assign decode_BYPASSABLE_MEMORY_STAGE = _zz_decode_IS_RS2_SIGNED[12];
  assign decode_BYPASSABLE_EXECUTE_STAGE = _zz_decode_IS_RS2_SIGNED[11];
  assign decode_SRC2_CTRL = _zz_decode_SRC2_CTRL;
  assign _zz_decode_to_execute_SRC2_CTRL = _zz_decode_to_execute_SRC2_CTRL_1;
  assign decode_ALU_CTRL = _zz_decode_ALU_CTRL;
  assign _zz_decode_to_execute_ALU_CTRL = _zz_decode_to_execute_ALU_CTRL_1;
  assign decode_SRC1_CTRL = _zz_decode_SRC1_CTRL;
  assign _zz_decode_to_execute_SRC1_CTRL = _zz_decode_to_execute_SRC1_CTRL_1;
  assign decode_MEMORY_FORCE_CONSTISTENCY = 1'b0;
  assign writeBack_FORMAL_PC_NEXT = memory_to_writeBack_FORMAL_PC_NEXT;
  assign memory_FORMAL_PC_NEXT = execute_to_memory_FORMAL_PC_NEXT;
  assign execute_FORMAL_PC_NEXT = decode_to_execute_FORMAL_PC_NEXT;
  assign decode_FORMAL_PC_NEXT = (decode_PC + 32'h00000004);
  assign memory_PC = execute_to_memory_PC;
  assign execute_IS_RS1_SIGNED = decode_to_execute_IS_RS1_SIGNED;
  assign execute_IS_DIV = decode_to_execute_IS_DIV;
  assign execute_IS_RS2_SIGNED = decode_to_execute_IS_RS2_SIGNED;
  assign memory_IS_DIV = execute_to_memory_IS_DIV;
  assign writeBack_IS_MUL = memory_to_writeBack_IS_MUL;
  assign writeBack_MUL_HH = memory_to_writeBack_MUL_HH;
  assign writeBack_MUL_LOW = memory_to_writeBack_MUL_LOW;
  assign memory_MUL_HL = execute_to_memory_MUL_HL;
  assign memory_MUL_LH = execute_to_memory_MUL_LH;
  assign memory_MUL_LL = execute_to_memory_MUL_LL;
  assign execute_CSR_READ_OPCODE = decode_to_execute_CSR_READ_OPCODE;
  assign execute_CSR_WRITE_OPCODE = decode_to_execute_CSR_WRITE_OPCODE;
  assign execute_IS_CSR = decode_to_execute_IS_CSR;
  assign memory_ENV_CTRL = _zz_memory_ENV_CTRL;
  assign execute_ENV_CTRL = _zz_execute_ENV_CTRL;
  assign writeBack_ENV_CTRL = _zz_writeBack_ENV_CTRL;
  assign memory_BRANCH_CALC = execute_to_memory_BRANCH_CALC;
  assign memory_BRANCH_DO = execute_to_memory_BRANCH_DO;
  assign execute_PC = decode_to_execute_PC;
  assign execute_PREDICTION_HAD_BRANCHED2 = decode_to_execute_PREDICTION_HAD_BRANCHED2;
  assign execute_BRANCH_COND_RESULT = _zz_execute_BRANCH_COND_RESULT_1;
  assign execute_BRANCH_CTRL = _zz_execute_BRANCH_CTRL;
  assign decode_RS2_USE = _zz_decode_IS_RS2_SIGNED[15];
  assign decode_RS1_USE = _zz_decode_IS_RS2_SIGNED[5];
  always @(*) begin
    _zz_decode_RS2 = execute_REGFILE_WRITE_DATA;
    if(when_CsrPlugin_l1189) begin
      _zz_decode_RS2 = CsrPlugin_csrMapping_readDataSignal;
    end
  end

  assign execute_REGFILE_WRITE_VALID = decode_to_execute_REGFILE_WRITE_VALID;
  assign execute_BYPASSABLE_EXECUTE_STAGE = decode_to_execute_BYPASSABLE_EXECUTE_STAGE;
  assign memory_REGFILE_WRITE_VALID = execute_to_memory_REGFILE_WRITE_VALID;
  assign memory_INSTRUCTION = execute_to_memory_INSTRUCTION;
  assign memory_BYPASSABLE_MEMORY_STAGE = execute_to_memory_BYPASSABLE_MEMORY_STAGE;
  assign writeBack_REGFILE_WRITE_VALID = memory_to_writeBack_REGFILE_WRITE_VALID;
  always @(*) begin
    decode_RS2 = decode_RegFilePlugin_rs2Data;
    if(HazardSimplePlugin_writeBackBuffer_valid) begin
      if(HazardSimplePlugin_addr1Match) begin
        decode_RS2 = HazardSimplePlugin_writeBackBuffer_payload_data;
      end
    end
    if(when_HazardSimplePlugin_l45) begin
      if(when_HazardSimplePlugin_l47) begin
        if(when_HazardSimplePlugin_l51) begin
          decode_RS2 = _zz_decode_RS2_2;
        end
      end
    end
    if(when_HazardSimplePlugin_l45_1) begin
      if(memory_BYPASSABLE_MEMORY_STAGE) begin
        if(when_HazardSimplePlugin_l51_1) begin
          decode_RS2 = _zz_decode_RS2_1;
        end
      end
    end
    if(when_HazardSimplePlugin_l45_2) begin
      if(execute_BYPASSABLE_EXECUTE_STAGE) begin
        if(when_HazardSimplePlugin_l51_2) begin
          decode_RS2 = _zz_decode_RS2;
        end
      end
    end
  end

  always @(*) begin
    decode_RS1 = decode_RegFilePlugin_rs1Data;
    if(HazardSimplePlugin_writeBackBuffer_valid) begin
      if(HazardSimplePlugin_addr0Match) begin
        decode_RS1 = HazardSimplePlugin_writeBackBuffer_payload_data;
      end
    end
    if(when_HazardSimplePlugin_l45) begin
      if(when_HazardSimplePlugin_l47) begin
        if(when_HazardSimplePlugin_l48) begin
          decode_RS1 = _zz_decode_RS2_2;
        end
      end
    end
    if(when_HazardSimplePlugin_l45_1) begin
      if(memory_BYPASSABLE_MEMORY_STAGE) begin
        if(when_HazardSimplePlugin_l48_1) begin
          decode_RS1 = _zz_decode_RS2_1;
        end
      end
    end
    if(when_HazardSimplePlugin_l45_2) begin
      if(execute_BYPASSABLE_EXECUTE_STAGE) begin
        if(when_HazardSimplePlugin_l48_2) begin
          decode_RS1 = _zz_decode_RS2;
        end
      end
    end
  end

  assign memory_SHIFT_RIGHT = execute_to_memory_SHIFT_RIGHT;
  always @(*) begin
    _zz_decode_RS2_1 = memory_REGFILE_WRITE_DATA;
    if(memory_arbitration_isValid) begin
      case(memory_SHIFT_CTRL)
        ShiftCtrlEnum_SLL_1 : begin
          _zz_decode_RS2_1 = _zz_decode_RS2_3;
        end
        ShiftCtrlEnum_SRL_1, ShiftCtrlEnum_SRA_1 : begin
          _zz_decode_RS2_1 = memory_SHIFT_RIGHT;
        end
        default : begin
        end
      endcase
    end
    if(when_MulDivIterativePlugin_l128) begin
      _zz_decode_RS2_1 = memory_DivPlugin_div_result;
    end
  end

  assign memory_SHIFT_CTRL = _zz_memory_SHIFT_CTRL;
  assign execute_SHIFT_CTRL = _zz_execute_SHIFT_CTRL;
  assign execute_SRC_LESS_UNSIGNED = decode_to_execute_SRC_LESS_UNSIGNED;
  assign execute_SRC2_FORCE_ZERO = decode_to_execute_SRC2_FORCE_ZERO;
  assign execute_SRC_USE_SUB_LESS = decode_to_execute_SRC_USE_SUB_LESS;
  assign _zz_execute_SRC2 = execute_PC;
  assign execute_SRC2_CTRL = _zz_execute_SRC2_CTRL;
  assign execute_SRC1_CTRL = _zz_execute_SRC1_CTRL;
  assign decode_SRC_USE_SUB_LESS = _zz_decode_IS_RS2_SIGNED[3];
  assign decode_SRC_ADD_ZERO = _zz_decode_IS_RS2_SIGNED[20];
  assign execute_SRC_ADD_SUB = execute_SrcPlugin_addSub;
  assign execute_SRC_LESS = execute_SrcPlugin_less;
  assign execute_ALU_CTRL = _zz_execute_ALU_CTRL;
  assign execute_SRC2 = _zz_execute_SRC2_5;
  assign execute_SRC1 = _zz_execute_SRC1;
  assign execute_ALU_BITWISE_CTRL = _zz_execute_ALU_BITWISE_CTRL;
  assign _zz_lastStageRegFileWrite_payload_address = writeBack_INSTRUCTION;
  assign _zz_lastStageRegFileWrite_valid = writeBack_REGFILE_WRITE_VALID;
  always @(*) begin
    _zz_2 = 1'b0;
    if(lastStageRegFileWrite_valid) begin
      _zz_2 = 1'b1;
    end
  end

  assign decode_INSTRUCTION_ANTICIPATED = (decode_arbitration_isStuck ? decode_INSTRUCTION : IBusCachedPlugin_cache_io_cpu_fetch_data);
  always @(*) begin
    decode_REGFILE_WRITE_VALID = _zz_decode_IS_RS2_SIGNED[10];
    if(when_RegFilePlugin_l63) begin
      decode_REGFILE_WRITE_VALID = 1'b0;
    end
  end

  assign decode_LEGAL_INSTRUCTION = (|{((decode_INSTRUCTION & 32'h0000005f) == 32'h00000017),{((decode_INSTRUCTION & 32'h0000007f) == 32'h0000006f),{((decode_INSTRUCTION & 32'h0000106f) == 32'h00000003),{((decode_INSTRUCTION & _zz_decode_LEGAL_INSTRUCTION) == 32'h00001073),{(_zz_decode_LEGAL_INSTRUCTION_1 == _zz_decode_LEGAL_INSTRUCTION_2),{_zz_decode_LEGAL_INSTRUCTION_3,{_zz_decode_LEGAL_INSTRUCTION_4,_zz_decode_LEGAL_INSTRUCTION_5}}}}}}});
  always @(*) begin
    _zz_decode_RS2_2 = writeBack_REGFILE_WRITE_DATA;
    if(when_DBusCachedPlugin_l492) begin
      _zz_decode_RS2_2 = writeBack_DBusCachedPlugin_rspFormated;
    end
    if(when_MulPlugin_l147) begin
      case(switch_MulPlugin_l148)
        2'b00 : begin
          _zz_decode_RS2_2 = _zz__zz_decode_RS2_2;
        end
        default : begin
          _zz_decode_RS2_2 = _zz__zz_decode_RS2_2_1;
        end
      endcase
    end
  end

  assign writeBack_MEMORY_WR = memory_to_writeBack_MEMORY_WR;
  assign writeBack_MEMORY_STORE_DATA_RF = memory_to_writeBack_MEMORY_STORE_DATA_RF;
  assign writeBack_REGFILE_WRITE_DATA = memory_to_writeBack_REGFILE_WRITE_DATA;
  assign writeBack_MEMORY_ENABLE = memory_to_writeBack_MEMORY_ENABLE;
  assign memory_REGFILE_WRITE_DATA = execute_to_memory_REGFILE_WRITE_DATA;
  assign memory_MEMORY_ENABLE = execute_to_memory_MEMORY_ENABLE;
  assign execute_MEMORY_FORCE_CONSTISTENCY = decode_to_execute_MEMORY_FORCE_CONSTISTENCY;
  assign execute_RS1 = decode_to_execute_RS1;
  assign execute_MEMORY_MANAGMENT = decode_to_execute_MEMORY_MANAGMENT;
  assign execute_RS2 = decode_to_execute_RS2;
  assign execute_MEMORY_WR = decode_to_execute_MEMORY_WR;
  assign execute_SRC_ADD = execute_SrcPlugin_addSub;
  assign execute_MEMORY_ENABLE = decode_to_execute_MEMORY_ENABLE;
  assign execute_INSTRUCTION = decode_to_execute_INSTRUCTION;
  assign decode_MEMORY_ENABLE = _zz_decode_IS_RS2_SIGNED[4];
  assign decode_FLUSH_ALL = _zz_decode_IS_RS2_SIGNED[0];
  always @(*) begin
    IBusCachedPlugin_rsp_issueDetected_4 = IBusCachedPlugin_rsp_issueDetected_3;
    if(when_IBusCachedPlugin_l256) begin
      IBusCachedPlugin_rsp_issueDetected_4 = 1'b1;
    end
  end

  always @(*) begin
    IBusCachedPlugin_rsp_issueDetected_3 = IBusCachedPlugin_rsp_issueDetected_2;
    if(when_IBusCachedPlugin_l250) begin
      IBusCachedPlugin_rsp_issueDetected_3 = 1'b1;
    end
  end

  always @(*) begin
    IBusCachedPlugin_rsp_issueDetected_2 = IBusCachedPlugin_rsp_issueDetected_1;
    if(when_IBusCachedPlugin_l244) begin
      IBusCachedPlugin_rsp_issueDetected_2 = 1'b1;
    end
  end

  always @(*) begin
    IBusCachedPlugin_rsp_issueDetected_1 = IBusCachedPlugin_rsp_issueDetected;
    if(when_IBusCachedPlugin_l239) begin
      IBusCachedPlugin_rsp_issueDetected_1 = 1'b1;
    end
  end

  assign decode_BRANCH_CTRL = _zz_decode_BRANCH_CTRL_1;
  assign decode_INSTRUCTION = IBusCachedPlugin_iBusRsp_output_payload_rsp_inst;
  always @(*) begin
    _zz_memory_to_writeBack_FORMAL_PC_NEXT = memory_FORMAL_PC_NEXT;
    if(BranchPlugin_jumpInterface_valid) begin
      _zz_memory_to_writeBack_FORMAL_PC_NEXT = BranchPlugin_jumpInterface_payload;
    end
  end

  always @(*) begin
    _zz_decode_to_execute_FORMAL_PC_NEXT = decode_FORMAL_PC_NEXT;
    if(IBusCachedPlugin_predictionJumpInterface_valid) begin
      _zz_decode_to_execute_FORMAL_PC_NEXT = IBusCachedPlugin_predictionJumpInterface_payload;
    end
  end

  assign decode_PC = IBusCachedPlugin_iBusRsp_output_payload_pc;
  assign writeBack_PC = memory_to_writeBack_PC;
  assign writeBack_INSTRUCTION = memory_to_writeBack_INSTRUCTION;
  always @(*) begin
    decode_arbitration_haltItself = 1'b0;
    if(when_DBusCachedPlugin_l308) begin
      decode_arbitration_haltItself = 1'b1;
    end
  end

  always @(*) begin
    decode_arbitration_haltByOther = 1'b0;
    if(when_HazardSimplePlugin_l113) begin
      decode_arbitration_haltByOther = 1'b1;
    end
    if(CsrPlugin_pipelineLiberator_active) begin
      decode_arbitration_haltByOther = 1'b1;
    end
    if(when_CsrPlugin_l1129) begin
      decode_arbitration_haltByOther = 1'b1;
    end
  end

  always @(*) begin
    decode_arbitration_removeIt = 1'b0;
    if(_zz_when) begin
      decode_arbitration_removeIt = 1'b1;
    end
    if(decode_arbitration_isFlushed) begin
      decode_arbitration_removeIt = 1'b1;
    end
  end

  assign decode_arbitration_flushIt = 1'b0;
  always @(*) begin
    decode_arbitration_flushNext = 1'b0;
    if(IBusCachedPlugin_predictionJumpInterface_valid) begin
      decode_arbitration_flushNext = 1'b1;
    end
    if(_zz_when) begin
      decode_arbitration_flushNext = 1'b1;
    end
  end

  always @(*) begin
    execute_arbitration_haltItself = 1'b0;
    if(when_DBusCachedPlugin_l350) begin
      execute_arbitration_haltItself = 1'b1;
    end
    if(when_CsrPlugin_l1121) begin
      if(when_CsrPlugin_l1123) begin
        execute_arbitration_haltItself = 1'b1;
      end
    end
    if(when_CsrPlugin_l1193) begin
      if(execute_CsrPlugin_blockedBySideEffects) begin
        execute_arbitration_haltItself = 1'b1;
      end
    end
    if(execute_CsrPlugin_writeInstruction) begin
      if(when_PmpPlugin_l172) begin
        execute_arbitration_haltItself = (! execute_PmpPlugin_fsmComplete);
      end
    end
  end

  always @(*) begin
    execute_arbitration_haltByOther = 1'b0;
    if(when_DBusCachedPlugin_l366) begin
      execute_arbitration_haltByOther = 1'b1;
    end
  end

  always @(*) begin
    execute_arbitration_removeIt = 1'b0;
    if(CsrPlugin_selfException_valid) begin
      execute_arbitration_removeIt = 1'b1;
    end
    if(execute_arbitration_isFlushed) begin
      execute_arbitration_removeIt = 1'b1;
    end
  end

  assign execute_arbitration_flushIt = 1'b0;
  always @(*) begin
    execute_arbitration_flushNext = 1'b0;
    if(CsrPlugin_selfException_valid) begin
      execute_arbitration_flushNext = 1'b1;
    end
  end

  always @(*) begin
    memory_arbitration_haltItself = 1'b0;
    if(when_MulDivIterativePlugin_l128) begin
      if(when_MulDivIterativePlugin_l129) begin
        memory_arbitration_haltItself = 1'b1;
      end
    end
  end

  assign memory_arbitration_haltByOther = 1'b0;
  always @(*) begin
    memory_arbitration_removeIt = 1'b0;
    if(BranchPlugin_branchExceptionPort_valid) begin
      memory_arbitration_removeIt = 1'b1;
    end
    if(memory_arbitration_isFlushed) begin
      memory_arbitration_removeIt = 1'b1;
    end
  end

  assign memory_arbitration_flushIt = 1'b0;
  always @(*) begin
    memory_arbitration_flushNext = 1'b0;
    if(BranchPlugin_jumpInterface_valid) begin
      memory_arbitration_flushNext = 1'b1;
    end
    if(BranchPlugin_branchExceptionPort_valid) begin
      memory_arbitration_flushNext = 1'b1;
    end
  end

  always @(*) begin
    writeBack_arbitration_haltItself = 1'b0;
    if(when_DBusCachedPlugin_l466) begin
      writeBack_arbitration_haltItself = 1'b1;
    end
  end

  assign writeBack_arbitration_haltByOther = 1'b0;
  always @(*) begin
    writeBack_arbitration_removeIt = 1'b0;
    if(DBusCachedPlugin_exceptionBus_valid) begin
      writeBack_arbitration_removeIt = 1'b1;
    end
    if(writeBack_arbitration_isFlushed) begin
      writeBack_arbitration_removeIt = 1'b1;
    end
  end

  always @(*) begin
    writeBack_arbitration_flushIt = 1'b0;
    if(DBusCachedPlugin_redoBranch_valid) begin
      writeBack_arbitration_flushIt = 1'b1;
    end
  end

  always @(*) begin
    writeBack_arbitration_flushNext = 1'b0;
    if(DBusCachedPlugin_redoBranch_valid) begin
      writeBack_arbitration_flushNext = 1'b1;
    end
    if(DBusCachedPlugin_exceptionBus_valid) begin
      writeBack_arbitration_flushNext = 1'b1;
    end
    if(when_CsrPlugin_l1032) begin
      writeBack_arbitration_flushNext = 1'b1;
    end
    if(when_CsrPlugin_l1077) begin
      writeBack_arbitration_flushNext = 1'b1;
    end
  end

  assign lastStageInstruction = writeBack_INSTRUCTION;
  assign lastStagePc = writeBack_PC;
  assign lastStageIsValid = writeBack_arbitration_isValid;
  assign lastStageIsFiring = writeBack_arbitration_isFiring;
  always @(*) begin
    IBusCachedPlugin_fetcherHalt = 1'b0;
    if(when_CsrPlugin_l935) begin
      IBusCachedPlugin_fetcherHalt = 1'b1;
    end
    if(when_CsrPlugin_l1032) begin
      IBusCachedPlugin_fetcherHalt = 1'b1;
    end
    if(when_CsrPlugin_l1077) begin
      IBusCachedPlugin_fetcherHalt = 1'b1;
    end
  end

  assign IBusCachedPlugin_forceNoDecodeCond = 1'b0;
  always @(*) begin
    IBusCachedPlugin_incomingInstruction = 1'b0;
    if(when_Fetcher_l243) begin
      IBusCachedPlugin_incomingInstruction = 1'b1;
    end
  end

  assign BranchPlugin_inDebugNoFetchFlag = 1'b0;
  always @(*) begin
    CsrPlugin_csrMapping_allowCsrSignal = 1'b0;
    if(execute_CsrPlugin_readInstruction) begin
      if(when_PmpPlugin_l155) begin
        if(execute_PmpPlugin_pmpcfgCsr) begin
          CsrPlugin_csrMapping_allowCsrSignal = 1'b1;
        end
        if(execute_PmpPlugin_pmpaddrCsr) begin
          CsrPlugin_csrMapping_allowCsrSignal = 1'b1;
        end
      end
    end
    if(execute_CsrPlugin_writeInstruction) begin
      if(when_PmpPlugin_l172) begin
        CsrPlugin_csrMapping_allowCsrSignal = 1'b1;
      end
    end
  end

  always @(*) begin
    CsrPlugin_csrMapping_readDataSignal = CsrPlugin_csrMapping_readDataInit;
    if(execute_CsrPlugin_readInstruction) begin
      if(when_PmpPlugin_l155) begin
        if(execute_PmpPlugin_pmpcfgCsr) begin
          CsrPlugin_csrMapping_readDataSignal = {{{_zz_CsrPlugin_csrMapping_readDataSignal,_zz_CsrPlugin_csrMapping_readDataSignal_2},_zz_CsrPlugin_csrMapping_readDataSignal_4},_zz_CsrPlugin_csrMapping_readDataSignal_6};
        end
        if(execute_PmpPlugin_pmpaddrCsr) begin
          CsrPlugin_csrMapping_readDataSignal = _zz_PmpPlugin_pmpaddr_port2;
        end
      end
    end
  end

  always @(*) begin
    CsrPlugin_inWfi = 1'b0;
    if(when_CsrPlugin_l1121) begin
      CsrPlugin_inWfi = 1'b1;
    end
  end

  assign CsrPlugin_thirdPartyWake = 1'b0;
  always @(*) begin
    CsrPlugin_jumpInterface_valid = 1'b0;
    if(when_CsrPlugin_l1032) begin
      CsrPlugin_jumpInterface_valid = 1'b1;
    end
    if(when_CsrPlugin_l1077) begin
      CsrPlugin_jumpInterface_valid = 1'b1;
    end
  end

  always @(*) begin
    CsrPlugin_jumpInterface_payload = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
    if(when_CsrPlugin_l1032) begin
      CsrPlugin_jumpInterface_payload = {CsrPlugin_xtvec_base,2'b00};
    end
    if(when_CsrPlugin_l1077) begin
      case(switch_CsrPlugin_l1081)
        2'b11 : begin
          CsrPlugin_jumpInterface_payload = CsrPlugin_mepc;
        end
        default : begin
        end
      endcase
    end
  end

  assign CsrPlugin_forceMachineWire = 1'b0;
  assign CsrPlugin_allowInterrupts = 1'b1;
  assign CsrPlugin_allowException = 1'b1;
  assign CsrPlugin_allowEbreakException = 1'b1;
  assign IBusCachedPlugin_externalFlush = ({writeBack_arbitration_flushNext,{memory_arbitration_flushNext,{execute_arbitration_flushNext,decode_arbitration_flushNext}}} != 4'b0000);
  assign IBusCachedPlugin_jump_pcLoad_valid = ({CsrPlugin_jumpInterface_valid,{BranchPlugin_jumpInterface_valid,{DBusCachedPlugin_redoBranch_valid,IBusCachedPlugin_predictionJumpInterface_valid}}} != 4'b0000);
  assign _zz_IBusCachedPlugin_jump_pcLoad_payload = {IBusCachedPlugin_predictionJumpInterface_valid,{BranchPlugin_jumpInterface_valid,{CsrPlugin_jumpInterface_valid,DBusCachedPlugin_redoBranch_valid}}};
  assign _zz_IBusCachedPlugin_jump_pcLoad_payload_1 = (_zz_IBusCachedPlugin_jump_pcLoad_payload & (~ _zz__zz_IBusCachedPlugin_jump_pcLoad_payload_1));
  assign _zz_IBusCachedPlugin_jump_pcLoad_payload_2 = _zz_IBusCachedPlugin_jump_pcLoad_payload_1[3];
  assign _zz_IBusCachedPlugin_jump_pcLoad_payload_3 = (_zz_IBusCachedPlugin_jump_pcLoad_payload_1[1] || _zz_IBusCachedPlugin_jump_pcLoad_payload_2);
  assign _zz_IBusCachedPlugin_jump_pcLoad_payload_4 = (_zz_IBusCachedPlugin_jump_pcLoad_payload_1[2] || _zz_IBusCachedPlugin_jump_pcLoad_payload_2);
  assign IBusCachedPlugin_jump_pcLoad_payload = _zz_IBusCachedPlugin_jump_pcLoad_payload_5;
  always @(*) begin
    IBusCachedPlugin_fetchPc_correction = 1'b0;
    if(IBusCachedPlugin_fetchPc_redo_valid) begin
      IBusCachedPlugin_fetchPc_correction = 1'b1;
    end
    if(IBusCachedPlugin_jump_pcLoad_valid) begin
      IBusCachedPlugin_fetchPc_correction = 1'b1;
    end
  end

  assign IBusCachedPlugin_fetchPc_output_fire = (IBusCachedPlugin_fetchPc_output_valid && IBusCachedPlugin_fetchPc_output_ready);
  assign IBusCachedPlugin_fetchPc_corrected = (IBusCachedPlugin_fetchPc_correction || IBusCachedPlugin_fetchPc_correctionReg);
  always @(*) begin
    IBusCachedPlugin_fetchPc_pcRegPropagate = 1'b0;
    if(IBusCachedPlugin_iBusRsp_stages_1_input_ready) begin
      IBusCachedPlugin_fetchPc_pcRegPropagate = 1'b1;
    end
  end

  assign when_Fetcher_l134 = (IBusCachedPlugin_fetchPc_correction || IBusCachedPlugin_fetchPc_pcRegPropagate);
  assign IBusCachedPlugin_fetchPc_output_fire_1 = (IBusCachedPlugin_fetchPc_output_valid && IBusCachedPlugin_fetchPc_output_ready);
  assign when_Fetcher_l134_1 = ((! IBusCachedPlugin_fetchPc_output_valid) && IBusCachedPlugin_fetchPc_output_ready);
  always @(*) begin
    IBusCachedPlugin_fetchPc_pc = (IBusCachedPlugin_fetchPc_pcReg + _zz_IBusCachedPlugin_fetchPc_pc);
    if(IBusCachedPlugin_fetchPc_redo_valid) begin
      IBusCachedPlugin_fetchPc_pc = IBusCachedPlugin_fetchPc_redo_payload;
    end
    if(IBusCachedPlugin_jump_pcLoad_valid) begin
      IBusCachedPlugin_fetchPc_pc = IBusCachedPlugin_jump_pcLoad_payload;
    end
    IBusCachedPlugin_fetchPc_pc[0] = 1'b0;
    IBusCachedPlugin_fetchPc_pc[1] = 1'b0;
  end

  always @(*) begin
    IBusCachedPlugin_fetchPc_flushed = 1'b0;
    if(IBusCachedPlugin_fetchPc_redo_valid) begin
      IBusCachedPlugin_fetchPc_flushed = 1'b1;
    end
    if(IBusCachedPlugin_jump_pcLoad_valid) begin
      IBusCachedPlugin_fetchPc_flushed = 1'b1;
    end
  end

  assign when_Fetcher_l161 = (IBusCachedPlugin_fetchPc_booted && ((IBusCachedPlugin_fetchPc_output_ready || IBusCachedPlugin_fetchPc_correction) || IBusCachedPlugin_fetchPc_pcRegPropagate));
  assign IBusCachedPlugin_fetchPc_output_valid = ((! IBusCachedPlugin_fetcherHalt) && IBusCachedPlugin_fetchPc_booted);
  assign IBusCachedPlugin_fetchPc_output_payload = IBusCachedPlugin_fetchPc_pc;
  always @(*) begin
    IBusCachedPlugin_iBusRsp_redoFetch = 1'b0;
    if(IBusCachedPlugin_rsp_redoFetch) begin
      IBusCachedPlugin_iBusRsp_redoFetch = 1'b1;
    end
  end

  assign IBusCachedPlugin_iBusRsp_stages_0_input_valid = IBusCachedPlugin_fetchPc_output_valid;
  assign IBusCachedPlugin_fetchPc_output_ready = IBusCachedPlugin_iBusRsp_stages_0_input_ready;
  assign IBusCachedPlugin_iBusRsp_stages_0_input_payload = IBusCachedPlugin_fetchPc_output_payload;
  always @(*) begin
    IBusCachedPlugin_iBusRsp_stages_0_halt = 1'b0;
    if(IBusCachedPlugin_cache_io_cpu_prefetch_haltIt) begin
      IBusCachedPlugin_iBusRsp_stages_0_halt = 1'b1;
    end
  end

  assign _zz_IBusCachedPlugin_iBusRsp_stages_0_input_ready = (! IBusCachedPlugin_iBusRsp_stages_0_halt);
  assign IBusCachedPlugin_iBusRsp_stages_0_input_ready = (IBusCachedPlugin_iBusRsp_stages_0_output_ready && _zz_IBusCachedPlugin_iBusRsp_stages_0_input_ready);
  assign IBusCachedPlugin_iBusRsp_stages_0_output_valid = (IBusCachedPlugin_iBusRsp_stages_0_input_valid && _zz_IBusCachedPlugin_iBusRsp_stages_0_input_ready);
  assign IBusCachedPlugin_iBusRsp_stages_0_output_payload = IBusCachedPlugin_iBusRsp_stages_0_input_payload;
  always @(*) begin
    IBusCachedPlugin_iBusRsp_stages_1_halt = 1'b0;
    if(IBusCachedPlugin_mmuBus_busy) begin
      IBusCachedPlugin_iBusRsp_stages_1_halt = 1'b1;
    end
  end

  assign _zz_IBusCachedPlugin_iBusRsp_stages_1_input_ready = (! IBusCachedPlugin_iBusRsp_stages_1_halt);
  assign IBusCachedPlugin_iBusRsp_stages_1_input_ready = (IBusCachedPlugin_iBusRsp_stages_1_output_ready && _zz_IBusCachedPlugin_iBusRsp_stages_1_input_ready);
  assign IBusCachedPlugin_iBusRsp_stages_1_output_valid = (IBusCachedPlugin_iBusRsp_stages_1_input_valid && _zz_IBusCachedPlugin_iBusRsp_stages_1_input_ready);
  assign IBusCachedPlugin_iBusRsp_stages_1_output_payload = IBusCachedPlugin_iBusRsp_stages_1_input_payload;
  always @(*) begin
    IBusCachedPlugin_iBusRsp_stages_2_halt = 1'b0;
    if(when_IBusCachedPlugin_l267) begin
      IBusCachedPlugin_iBusRsp_stages_2_halt = 1'b1;
    end
  end

  assign _zz_IBusCachedPlugin_iBusRsp_stages_2_input_ready = (! IBusCachedPlugin_iBusRsp_stages_2_halt);
  assign IBusCachedPlugin_iBusRsp_stages_2_input_ready = (IBusCachedPlugin_iBusRsp_stages_2_output_ready && _zz_IBusCachedPlugin_iBusRsp_stages_2_input_ready);
  assign IBusCachedPlugin_iBusRsp_stages_2_output_valid = (IBusCachedPlugin_iBusRsp_stages_2_input_valid && _zz_IBusCachedPlugin_iBusRsp_stages_2_input_ready);
  assign IBusCachedPlugin_iBusRsp_stages_2_output_payload = IBusCachedPlugin_iBusRsp_stages_2_input_payload;
  assign IBusCachedPlugin_fetchPc_redo_valid = IBusCachedPlugin_iBusRsp_redoFetch;
  assign IBusCachedPlugin_fetchPc_redo_payload = IBusCachedPlugin_iBusRsp_stages_2_input_payload;
  assign IBusCachedPlugin_iBusRsp_flush = ((decode_arbitration_removeIt || (decode_arbitration_flushNext && (! decode_arbitration_isStuck))) || IBusCachedPlugin_iBusRsp_redoFetch);
  assign IBusCachedPlugin_iBusRsp_stages_0_output_ready = _zz_IBusCachedPlugin_iBusRsp_stages_0_output_ready;
  assign _zz_IBusCachedPlugin_iBusRsp_stages_0_output_ready = ((1'b0 && (! _zz_IBusCachedPlugin_iBusRsp_stages_0_output_ready_1)) || IBusCachedPlugin_iBusRsp_stages_1_input_ready);
  assign _zz_IBusCachedPlugin_iBusRsp_stages_0_output_ready_1 = _zz_IBusCachedPlugin_iBusRsp_stages_0_output_ready_2;
  assign IBusCachedPlugin_iBusRsp_stages_1_input_valid = _zz_IBusCachedPlugin_iBusRsp_stages_0_output_ready_1;
  assign IBusCachedPlugin_iBusRsp_stages_1_input_payload = IBusCachedPlugin_fetchPc_pcReg;
  assign IBusCachedPlugin_iBusRsp_stages_1_output_ready = ((1'b0 && (! IBusCachedPlugin_iBusRsp_stages_1_output_m2sPipe_valid)) || IBusCachedPlugin_iBusRsp_stages_1_output_m2sPipe_ready);
  assign IBusCachedPlugin_iBusRsp_stages_1_output_m2sPipe_valid = _zz_IBusCachedPlugin_iBusRsp_stages_1_output_m2sPipe_valid;
  assign IBusCachedPlugin_iBusRsp_stages_1_output_m2sPipe_payload = _zz_IBusCachedPlugin_iBusRsp_stages_1_output_m2sPipe_payload;
  assign IBusCachedPlugin_iBusRsp_stages_2_input_valid = IBusCachedPlugin_iBusRsp_stages_1_output_m2sPipe_valid;
  assign IBusCachedPlugin_iBusRsp_stages_1_output_m2sPipe_ready = IBusCachedPlugin_iBusRsp_stages_2_input_ready;
  assign IBusCachedPlugin_iBusRsp_stages_2_input_payload = IBusCachedPlugin_iBusRsp_stages_1_output_m2sPipe_payload;
  always @(*) begin
    IBusCachedPlugin_iBusRsp_readyForError = 1'b1;
    if(when_Fetcher_l323) begin
      IBusCachedPlugin_iBusRsp_readyForError = 1'b0;
    end
  end

  assign when_Fetcher_l243 = (IBusCachedPlugin_iBusRsp_stages_1_input_valid || IBusCachedPlugin_iBusRsp_stages_2_input_valid);
  assign when_Fetcher_l323 = (! IBusCachedPlugin_pcValids_0);
  assign when_Fetcher_l332 = (! (! IBusCachedPlugin_iBusRsp_stages_1_input_ready));
  assign when_Fetcher_l332_1 = (! (! IBusCachedPlugin_iBusRsp_stages_2_input_ready));
  assign when_Fetcher_l332_2 = (! execute_arbitration_isStuck);
  assign when_Fetcher_l332_3 = (! memory_arbitration_isStuck);
  assign when_Fetcher_l332_4 = (! writeBack_arbitration_isStuck);
  assign IBusCachedPlugin_pcValids_0 = IBusCachedPlugin_injector_nextPcCalc_valids_1;
  assign IBusCachedPlugin_pcValids_1 = IBusCachedPlugin_injector_nextPcCalc_valids_2;
  assign IBusCachedPlugin_pcValids_2 = IBusCachedPlugin_injector_nextPcCalc_valids_3;
  assign IBusCachedPlugin_pcValids_3 = IBusCachedPlugin_injector_nextPcCalc_valids_4;
  assign IBusCachedPlugin_iBusRsp_output_ready = (! decode_arbitration_isStuck);
  always @(*) begin
    decode_arbitration_isValid = IBusCachedPlugin_iBusRsp_output_valid;
    if(IBusCachedPlugin_forceNoDecodeCond) begin
      decode_arbitration_isValid = 1'b0;
    end
  end

  assign _zz_IBusCachedPlugin_decodePrediction_cmd_hadBranch = _zz__zz_IBusCachedPlugin_decodePrediction_cmd_hadBranch[11];
  always @(*) begin
    _zz_IBusCachedPlugin_decodePrediction_cmd_hadBranch_1[18] = _zz_IBusCachedPlugin_decodePrediction_cmd_hadBranch;
    _zz_IBusCachedPlugin_decodePrediction_cmd_hadBranch_1[17] = _zz_IBusCachedPlugin_decodePrediction_cmd_hadBranch;
    _zz_IBusCachedPlugin_decodePrediction_cmd_hadBranch_1[16] = _zz_IBusCachedPlugin_decodePrediction_cmd_hadBranch;
    _zz_IBusCachedPlugin_decodePrediction_cmd_hadBranch_1[15] = _zz_IBusCachedPlugin_decodePrediction_cmd_hadBranch;
    _zz_IBusCachedPlugin_decodePrediction_cmd_hadBranch_1[14] = _zz_IBusCachedPlugin_decodePrediction_cmd_hadBranch;
    _zz_IBusCachedPlugin_decodePrediction_cmd_hadBranch_1[13] = _zz_IBusCachedPlugin_decodePrediction_cmd_hadBranch;
    _zz_IBusCachedPlugin_decodePrediction_cmd_hadBranch_1[12] = _zz_IBusCachedPlugin_decodePrediction_cmd_hadBranch;
    _zz_IBusCachedPlugin_decodePrediction_cmd_hadBranch_1[11] = _zz_IBusCachedPlugin_decodePrediction_cmd_hadBranch;
    _zz_IBusCachedPlugin_decodePrediction_cmd_hadBranch_1[10] = _zz_IBusCachedPlugin_decodePrediction_cmd_hadBranch;
    _zz_IBusCachedPlugin_decodePrediction_cmd_hadBranch_1[9] = _zz_IBusCachedPlugin_decodePrediction_cmd_hadBranch;
    _zz_IBusCachedPlugin_decodePrediction_cmd_hadBranch_1[8] = _zz_IBusCachedPlugin_decodePrediction_cmd_hadBranch;
    _zz_IBusCachedPlugin_decodePrediction_cmd_hadBranch_1[7] = _zz_IBusCachedPlugin_decodePrediction_cmd_hadBranch;
    _zz_IBusCachedPlugin_decodePrediction_cmd_hadBranch_1[6] = _zz_IBusCachedPlugin_decodePrediction_cmd_hadBranch;
    _zz_IBusCachedPlugin_decodePrediction_cmd_hadBranch_1[5] = _zz_IBusCachedPlugin_decodePrediction_cmd_hadBranch;
    _zz_IBusCachedPlugin_decodePrediction_cmd_hadBranch_1[4] = _zz_IBusCachedPlugin_decodePrediction_cmd_hadBranch;
    _zz_IBusCachedPlugin_decodePrediction_cmd_hadBranch_1[3] = _zz_IBusCachedPlugin_decodePrediction_cmd_hadBranch;
    _zz_IBusCachedPlugin_decodePrediction_cmd_hadBranch_1[2] = _zz_IBusCachedPlugin_decodePrediction_cmd_hadBranch;
    _zz_IBusCachedPlugin_decodePrediction_cmd_hadBranch_1[1] = _zz_IBusCachedPlugin_decodePrediction_cmd_hadBranch;
    _zz_IBusCachedPlugin_decodePrediction_cmd_hadBranch_1[0] = _zz_IBusCachedPlugin_decodePrediction_cmd_hadBranch;
  end

  always @(*) begin
    IBusCachedPlugin_decodePrediction_cmd_hadBranch = ((decode_BRANCH_CTRL == BranchCtrlEnum_JAL) || ((decode_BRANCH_CTRL == BranchCtrlEnum_B) && _zz_IBusCachedPlugin_decodePrediction_cmd_hadBranch_2[31]));
    if(_zz_7) begin
      IBusCachedPlugin_decodePrediction_cmd_hadBranch = 1'b0;
    end
  end

  assign _zz_3 = _zz__zz_3[19];
  always @(*) begin
    _zz_4[10] = _zz_3;
    _zz_4[9] = _zz_3;
    _zz_4[8] = _zz_3;
    _zz_4[7] = _zz_3;
    _zz_4[6] = _zz_3;
    _zz_4[5] = _zz_3;
    _zz_4[4] = _zz_3;
    _zz_4[3] = _zz_3;
    _zz_4[2] = _zz_3;
    _zz_4[1] = _zz_3;
    _zz_4[0] = _zz_3;
  end

  assign _zz_5 = _zz__zz_5[11];
  always @(*) begin
    _zz_6[18] = _zz_5;
    _zz_6[17] = _zz_5;
    _zz_6[16] = _zz_5;
    _zz_6[15] = _zz_5;
    _zz_6[14] = _zz_5;
    _zz_6[13] = _zz_5;
    _zz_6[12] = _zz_5;
    _zz_6[11] = _zz_5;
    _zz_6[10] = _zz_5;
    _zz_6[9] = _zz_5;
    _zz_6[8] = _zz_5;
    _zz_6[7] = _zz_5;
    _zz_6[6] = _zz_5;
    _zz_6[5] = _zz_5;
    _zz_6[4] = _zz_5;
    _zz_6[3] = _zz_5;
    _zz_6[2] = _zz_5;
    _zz_6[1] = _zz_5;
    _zz_6[0] = _zz_5;
  end

  always @(*) begin
    case(decode_BRANCH_CTRL)
      BranchCtrlEnum_JAL : begin
        _zz_7 = _zz__zz_7[1];
      end
      default : begin
        _zz_7 = _zz__zz_7_1[1];
      end
    endcase
  end

  assign IBusCachedPlugin_predictionJumpInterface_valid = (decode_arbitration_isValid && IBusCachedPlugin_decodePrediction_cmd_hadBranch);
  assign _zz_IBusCachedPlugin_predictionJumpInterface_payload = _zz__zz_IBusCachedPlugin_predictionJumpInterface_payload[19];
  always @(*) begin
    _zz_IBusCachedPlugin_predictionJumpInterface_payload_1[10] = _zz_IBusCachedPlugin_predictionJumpInterface_payload;
    _zz_IBusCachedPlugin_predictionJumpInterface_payload_1[9] = _zz_IBusCachedPlugin_predictionJumpInterface_payload;
    _zz_IBusCachedPlugin_predictionJumpInterface_payload_1[8] = _zz_IBusCachedPlugin_predictionJumpInterface_payload;
    _zz_IBusCachedPlugin_predictionJumpInterface_payload_1[7] = _zz_IBusCachedPlugin_predictionJumpInterface_payload;
    _zz_IBusCachedPlugin_predictionJumpInterface_payload_1[6] = _zz_IBusCachedPlugin_predictionJumpInterface_payload;
    _zz_IBusCachedPlugin_predictionJumpInterface_payload_1[5] = _zz_IBusCachedPlugin_predictionJumpInterface_payload;
    _zz_IBusCachedPlugin_predictionJumpInterface_payload_1[4] = _zz_IBusCachedPlugin_predictionJumpInterface_payload;
    _zz_IBusCachedPlugin_predictionJumpInterface_payload_1[3] = _zz_IBusCachedPlugin_predictionJumpInterface_payload;
    _zz_IBusCachedPlugin_predictionJumpInterface_payload_1[2] = _zz_IBusCachedPlugin_predictionJumpInterface_payload;
    _zz_IBusCachedPlugin_predictionJumpInterface_payload_1[1] = _zz_IBusCachedPlugin_predictionJumpInterface_payload;
    _zz_IBusCachedPlugin_predictionJumpInterface_payload_1[0] = _zz_IBusCachedPlugin_predictionJumpInterface_payload;
  end

  assign _zz_IBusCachedPlugin_predictionJumpInterface_payload_2 = _zz__zz_IBusCachedPlugin_predictionJumpInterface_payload_2[11];
  always @(*) begin
    _zz_IBusCachedPlugin_predictionJumpInterface_payload_3[18] = _zz_IBusCachedPlugin_predictionJumpInterface_payload_2;
    _zz_IBusCachedPlugin_predictionJumpInterface_payload_3[17] = _zz_IBusCachedPlugin_predictionJumpInterface_payload_2;
    _zz_IBusCachedPlugin_predictionJumpInterface_payload_3[16] = _zz_IBusCachedPlugin_predictionJumpInterface_payload_2;
    _zz_IBusCachedPlugin_predictionJumpInterface_payload_3[15] = _zz_IBusCachedPlugin_predictionJumpInterface_payload_2;
    _zz_IBusCachedPlugin_predictionJumpInterface_payload_3[14] = _zz_IBusCachedPlugin_predictionJumpInterface_payload_2;
    _zz_IBusCachedPlugin_predictionJumpInterface_payload_3[13] = _zz_IBusCachedPlugin_predictionJumpInterface_payload_2;
    _zz_IBusCachedPlugin_predictionJumpInterface_payload_3[12] = _zz_IBusCachedPlugin_predictionJumpInterface_payload_2;
    _zz_IBusCachedPlugin_predictionJumpInterface_payload_3[11] = _zz_IBusCachedPlugin_predictionJumpInterface_payload_2;
    _zz_IBusCachedPlugin_predictionJumpInterface_payload_3[10] = _zz_IBusCachedPlugin_predictionJumpInterface_payload_2;
    _zz_IBusCachedPlugin_predictionJumpInterface_payload_3[9] = _zz_IBusCachedPlugin_predictionJumpInterface_payload_2;
    _zz_IBusCachedPlugin_predictionJumpInterface_payload_3[8] = _zz_IBusCachedPlugin_predictionJumpInterface_payload_2;
    _zz_IBusCachedPlugin_predictionJumpInterface_payload_3[7] = _zz_IBusCachedPlugin_predictionJumpInterface_payload_2;
    _zz_IBusCachedPlugin_predictionJumpInterface_payload_3[6] = _zz_IBusCachedPlugin_predictionJumpInterface_payload_2;
    _zz_IBusCachedPlugin_predictionJumpInterface_payload_3[5] = _zz_IBusCachedPlugin_predictionJumpInterface_payload_2;
    _zz_IBusCachedPlugin_predictionJumpInterface_payload_3[4] = _zz_IBusCachedPlugin_predictionJumpInterface_payload_2;
    _zz_IBusCachedPlugin_predictionJumpInterface_payload_3[3] = _zz_IBusCachedPlugin_predictionJumpInterface_payload_2;
    _zz_IBusCachedPlugin_predictionJumpInterface_payload_3[2] = _zz_IBusCachedPlugin_predictionJumpInterface_payload_2;
    _zz_IBusCachedPlugin_predictionJumpInterface_payload_3[1] = _zz_IBusCachedPlugin_predictionJumpInterface_payload_2;
    _zz_IBusCachedPlugin_predictionJumpInterface_payload_3[0] = _zz_IBusCachedPlugin_predictionJumpInterface_payload_2;
  end

  assign IBusCachedPlugin_predictionJumpInterface_payload = (decode_PC + ((decode_BRANCH_CTRL == BranchCtrlEnum_JAL) ? {{_zz_IBusCachedPlugin_predictionJumpInterface_payload_1,{{{_zz_IBusCachedPlugin_predictionJumpInterface_payload_4,decode_INSTRUCTION[19 : 12]},decode_INSTRUCTION[20]},decode_INSTRUCTION[30 : 21]}},1'b0} : {{_zz_IBusCachedPlugin_predictionJumpInterface_payload_3,{{{_zz_IBusCachedPlugin_predictionJumpInterface_payload_5,_zz_IBusCachedPlugin_predictionJumpInterface_payload_6},decode_INSTRUCTION[30 : 25]},decode_INSTRUCTION[11 : 8]}},1'b0}));
  assign iBus_cmd_valid = IBusCachedPlugin_cache_io_mem_cmd_valid;
  always @(*) begin
    iBus_cmd_payload_address = IBusCachedPlugin_cache_io_mem_cmd_payload_address;
    iBus_cmd_payload_address = IBusCachedPlugin_cache_io_mem_cmd_payload_address;
  end

  assign iBus_cmd_payload_size = IBusCachedPlugin_cache_io_mem_cmd_payload_size;
  assign IBusCachedPlugin_s0_tightlyCoupledHit = 1'b0;
  assign IBusCachedPlugin_cache_io_cpu_prefetch_isValid = (IBusCachedPlugin_iBusRsp_stages_0_input_valid && (! IBusCachedPlugin_s0_tightlyCoupledHit));
  assign IBusCachedPlugin_cache_io_cpu_fetch_isValid = (IBusCachedPlugin_iBusRsp_stages_1_input_valid && (! IBusCachedPlugin_s1_tightlyCoupledHit));
  assign IBusCachedPlugin_cache_io_cpu_fetch_isStuck = (! IBusCachedPlugin_iBusRsp_stages_1_input_ready);
  assign IBusCachedPlugin_mmuBus_cmd_0_isValid = IBusCachedPlugin_cache_io_cpu_fetch_isValid;
  assign IBusCachedPlugin_mmuBus_cmd_0_isStuck = (! IBusCachedPlugin_iBusRsp_stages_1_input_ready);
  assign IBusCachedPlugin_mmuBus_cmd_0_virtualAddress = IBusCachedPlugin_iBusRsp_stages_1_input_payload;
  assign IBusCachedPlugin_mmuBus_cmd_0_bypassTranslation = 1'b0;
  assign IBusCachedPlugin_mmuBus_end = (IBusCachedPlugin_iBusRsp_stages_1_input_ready || IBusCachedPlugin_externalFlush);
  assign IBusCachedPlugin_cache_io_cpu_decode_isValid = (IBusCachedPlugin_iBusRsp_stages_2_input_valid && (! IBusCachedPlugin_s2_tightlyCoupledHit));
  assign IBusCachedPlugin_cache_io_cpu_decode_isStuck = (! IBusCachedPlugin_iBusRsp_stages_2_input_ready);
  assign IBusCachedPlugin_cache_io_cpu_decode_isUser = (CsrPlugin_privilege == 2'b00);
  assign IBusCachedPlugin_rsp_iBusRspOutputHalt = 1'b0;
  assign IBusCachedPlugin_rsp_issueDetected = 1'b0;
  always @(*) begin
    IBusCachedPlugin_rsp_redoFetch = 1'b0;
    if(when_IBusCachedPlugin_l239) begin
      IBusCachedPlugin_rsp_redoFetch = 1'b1;
    end
    if(when_IBusCachedPlugin_l250) begin
      IBusCachedPlugin_rsp_redoFetch = 1'b1;
    end
  end

  always @(*) begin
    IBusCachedPlugin_cache_io_cpu_fill_valid = (IBusCachedPlugin_rsp_redoFetch && (! IBusCachedPlugin_cache_io_cpu_decode_mmuRefilling));
    if(when_IBusCachedPlugin_l250) begin
      IBusCachedPlugin_cache_io_cpu_fill_valid = 1'b1;
    end
  end

  always @(*) begin
    IBusCachedPlugin_decodeExceptionPort_valid = 1'b0;
    if(when_IBusCachedPlugin_l244) begin
      IBusCachedPlugin_decodeExceptionPort_valid = IBusCachedPlugin_iBusRsp_readyForError;
    end
    if(when_IBusCachedPlugin_l256) begin
      IBusCachedPlugin_decodeExceptionPort_valid = IBusCachedPlugin_iBusRsp_readyForError;
    end
  end

  always @(*) begin
    IBusCachedPlugin_decodeExceptionPort_payload_code = 4'bxxxx;
    if(when_IBusCachedPlugin_l244) begin
      IBusCachedPlugin_decodeExceptionPort_payload_code = 4'b1100;
    end
    if(when_IBusCachedPlugin_l256) begin
      IBusCachedPlugin_decodeExceptionPort_payload_code = 4'b0001;
    end
  end

  assign IBusCachedPlugin_decodeExceptionPort_payload_badAddr = {IBusCachedPlugin_iBusRsp_stages_2_input_payload[31 : 2],2'b00};
  assign when_IBusCachedPlugin_l239 = ((IBusCachedPlugin_cache_io_cpu_decode_isValid && IBusCachedPlugin_cache_io_cpu_decode_mmuRefilling) && (! IBusCachedPlugin_rsp_issueDetected));
  assign when_IBusCachedPlugin_l244 = ((IBusCachedPlugin_cache_io_cpu_decode_isValid && IBusCachedPlugin_cache_io_cpu_decode_mmuException) && (! IBusCachedPlugin_rsp_issueDetected_1));
  assign when_IBusCachedPlugin_l250 = ((IBusCachedPlugin_cache_io_cpu_decode_isValid && IBusCachedPlugin_cache_io_cpu_decode_cacheMiss) && (! IBusCachedPlugin_rsp_issueDetected_2));
  assign when_IBusCachedPlugin_l256 = ((IBusCachedPlugin_cache_io_cpu_decode_isValid && IBusCachedPlugin_cache_io_cpu_decode_error) && (! IBusCachedPlugin_rsp_issueDetected_3));
  assign when_IBusCachedPlugin_l267 = (IBusCachedPlugin_rsp_issueDetected_4 || IBusCachedPlugin_rsp_iBusRspOutputHalt);
  assign IBusCachedPlugin_iBusRsp_output_valid = IBusCachedPlugin_iBusRsp_stages_2_output_valid;
  assign IBusCachedPlugin_iBusRsp_stages_2_output_ready = IBusCachedPlugin_iBusRsp_output_ready;
  assign IBusCachedPlugin_iBusRsp_output_payload_rsp_inst = IBusCachedPlugin_cache_io_cpu_decode_data;
  assign IBusCachedPlugin_iBusRsp_output_payload_pc = IBusCachedPlugin_iBusRsp_stages_2_output_payload;
  assign IBusCachedPlugin_cache_io_flush = (decode_arbitration_isValid && decode_FLUSH_ALL);
  assign dataCache_1_io_mem_cmd_ready = (! dataCache_1_io_mem_cmd_rValid);
  assign dataCache_1_io_mem_cmd_s2mPipe_valid = (dataCache_1_io_mem_cmd_valid || dataCache_1_io_mem_cmd_rValid);
  assign dataCache_1_io_mem_cmd_s2mPipe_payload_wr = (dataCache_1_io_mem_cmd_rValid ? dataCache_1_io_mem_cmd_rData_wr : dataCache_1_io_mem_cmd_payload_wr);
  assign dataCache_1_io_mem_cmd_s2mPipe_payload_uncached = (dataCache_1_io_mem_cmd_rValid ? dataCache_1_io_mem_cmd_rData_uncached : dataCache_1_io_mem_cmd_payload_uncached);
  assign dataCache_1_io_mem_cmd_s2mPipe_payload_address = (dataCache_1_io_mem_cmd_rValid ? dataCache_1_io_mem_cmd_rData_address : dataCache_1_io_mem_cmd_payload_address);
  assign dataCache_1_io_mem_cmd_s2mPipe_payload_data = (dataCache_1_io_mem_cmd_rValid ? dataCache_1_io_mem_cmd_rData_data : dataCache_1_io_mem_cmd_payload_data);
  assign dataCache_1_io_mem_cmd_s2mPipe_payload_mask = (dataCache_1_io_mem_cmd_rValid ? dataCache_1_io_mem_cmd_rData_mask : dataCache_1_io_mem_cmd_payload_mask);
  assign dataCache_1_io_mem_cmd_s2mPipe_payload_size = (dataCache_1_io_mem_cmd_rValid ? dataCache_1_io_mem_cmd_rData_size : dataCache_1_io_mem_cmd_payload_size);
  assign dataCache_1_io_mem_cmd_s2mPipe_payload_last = (dataCache_1_io_mem_cmd_rValid ? dataCache_1_io_mem_cmd_rData_last : dataCache_1_io_mem_cmd_payload_last);
  always @(*) begin
    dataCache_1_io_mem_cmd_s2mPipe_ready = dataCache_1_io_mem_cmd_s2mPipe_m2sPipe_ready;
    if(when_Stream_l368) begin
      dataCache_1_io_mem_cmd_s2mPipe_ready = 1'b1;
    end
  end

  assign when_Stream_l368 = (! dataCache_1_io_mem_cmd_s2mPipe_m2sPipe_valid);
  assign dataCache_1_io_mem_cmd_s2mPipe_m2sPipe_valid = dataCache_1_io_mem_cmd_s2mPipe_rValid;
  assign dataCache_1_io_mem_cmd_s2mPipe_m2sPipe_payload_wr = dataCache_1_io_mem_cmd_s2mPipe_rData_wr;
  assign dataCache_1_io_mem_cmd_s2mPipe_m2sPipe_payload_uncached = dataCache_1_io_mem_cmd_s2mPipe_rData_uncached;
  assign dataCache_1_io_mem_cmd_s2mPipe_m2sPipe_payload_address = dataCache_1_io_mem_cmd_s2mPipe_rData_address;
  assign dataCache_1_io_mem_cmd_s2mPipe_m2sPipe_payload_data = dataCache_1_io_mem_cmd_s2mPipe_rData_data;
  assign dataCache_1_io_mem_cmd_s2mPipe_m2sPipe_payload_mask = dataCache_1_io_mem_cmd_s2mPipe_rData_mask;
  assign dataCache_1_io_mem_cmd_s2mPipe_m2sPipe_payload_size = dataCache_1_io_mem_cmd_s2mPipe_rData_size;
  assign dataCache_1_io_mem_cmd_s2mPipe_m2sPipe_payload_last = dataCache_1_io_mem_cmd_s2mPipe_rData_last;
  assign dBus_cmd_valid = dataCache_1_io_mem_cmd_s2mPipe_m2sPipe_valid;
  assign dataCache_1_io_mem_cmd_s2mPipe_m2sPipe_ready = dBus_cmd_ready;
  assign dBus_cmd_payload_wr = dataCache_1_io_mem_cmd_s2mPipe_m2sPipe_payload_wr;
  assign dBus_cmd_payload_uncached = dataCache_1_io_mem_cmd_s2mPipe_m2sPipe_payload_uncached;
  assign dBus_cmd_payload_address = dataCache_1_io_mem_cmd_s2mPipe_m2sPipe_payload_address;
  assign dBus_cmd_payload_data = dataCache_1_io_mem_cmd_s2mPipe_m2sPipe_payload_data;
  assign dBus_cmd_payload_mask = dataCache_1_io_mem_cmd_s2mPipe_m2sPipe_payload_mask;
  assign dBus_cmd_payload_size = dataCache_1_io_mem_cmd_s2mPipe_m2sPipe_payload_size;
  assign dBus_cmd_payload_last = dataCache_1_io_mem_cmd_s2mPipe_m2sPipe_payload_last;
  assign when_DBusCachedPlugin_l308 = ((DBusCachedPlugin_mmuBus_busy && decode_arbitration_isValid) && decode_MEMORY_ENABLE);
  assign execute_DBusCachedPlugin_size = execute_INSTRUCTION[13 : 12];
  assign dataCache_1_io_cpu_execute_isValid = (execute_arbitration_isValid && execute_MEMORY_ENABLE);
  assign dataCache_1_io_cpu_execute_address = execute_SRC_ADD;
  always @(*) begin
    case(execute_DBusCachedPlugin_size)
      2'b00 : begin
        _zz_execute_MEMORY_STORE_DATA_RF = {{{execute_RS2[7 : 0],execute_RS2[7 : 0]},execute_RS2[7 : 0]},execute_RS2[7 : 0]};
      end
      2'b01 : begin
        _zz_execute_MEMORY_STORE_DATA_RF = {execute_RS2[15 : 0],execute_RS2[15 : 0]};
      end
      default : begin
        _zz_execute_MEMORY_STORE_DATA_RF = execute_RS2[31 : 0];
      end
    endcase
  end

  assign dataCache_1_io_cpu_flush_valid = (execute_arbitration_isValid && execute_MEMORY_MANAGMENT);
  assign dataCache_1_io_cpu_flush_payload_singleLine = (execute_INSTRUCTION[19 : 15] != 5'h0);
  assign dataCache_1_io_cpu_flush_payload_lineId = _zz_io_cpu_flush_payload_lineId[6:0];
  assign dataCache_1_io_cpu_flush_isStall = (dataCache_1_io_cpu_flush_valid && (! dataCache_1_io_cpu_flush_ready));
  assign when_DBusCachedPlugin_l350 = (dataCache_1_io_cpu_flush_isStall || dataCache_1_io_cpu_execute_haltIt);
  assign when_DBusCachedPlugin_l366 = (dataCache_1_io_cpu_execute_refilling && execute_arbitration_isValid);
  assign dataCache_1_io_cpu_memory_isValid = (memory_arbitration_isValid && memory_MEMORY_ENABLE);
  assign dataCache_1_io_cpu_memory_address = memory_REGFILE_WRITE_DATA;
  assign DBusCachedPlugin_mmuBus_cmd_0_isValid = dataCache_1_io_cpu_memory_isValid;
  assign DBusCachedPlugin_mmuBus_cmd_0_isStuck = memory_arbitration_isStuck;
  assign DBusCachedPlugin_mmuBus_cmd_0_virtualAddress = dataCache_1_io_cpu_memory_address;
  assign DBusCachedPlugin_mmuBus_cmd_0_bypassTranslation = 1'b0;
  assign DBusCachedPlugin_mmuBus_end = ((! memory_arbitration_isStuck) || memory_arbitration_removeIt);
  always @(*) begin
    dataCache_1_io_cpu_memory_mmuRsp_isIoAccess = DBusCachedPlugin_mmuBus_rsp_isIoAccess;
    if(when_DBusCachedPlugin_l393) begin
      dataCache_1_io_cpu_memory_mmuRsp_isIoAccess = 1'b1;
    end
  end

  assign when_DBusCachedPlugin_l393 = (1'b0 && (! dataCache_1_io_cpu_memory_isWrite));
  always @(*) begin
    dataCache_1_io_cpu_writeBack_isValid = (writeBack_arbitration_isValid && writeBack_MEMORY_ENABLE);
    if(writeBack_arbitration_haltByOther) begin
      dataCache_1_io_cpu_writeBack_isValid = 1'b0;
    end
  end

  assign dataCache_1_io_cpu_writeBack_isUser = (CsrPlugin_privilege == 2'b00);
  assign dataCache_1_io_cpu_writeBack_address = writeBack_REGFILE_WRITE_DATA;
  assign dataCache_1_io_cpu_writeBack_storeData[31 : 0] = writeBack_MEMORY_STORE_DATA_RF;
  always @(*) begin
    DBusCachedPlugin_redoBranch_valid = 1'b0;
    if(when_DBusCachedPlugin_l446) begin
      if(dataCache_1_io_cpu_redo) begin
        DBusCachedPlugin_redoBranch_valid = 1'b1;
      end
    end
  end

  assign DBusCachedPlugin_redoBranch_payload = writeBack_PC;
  always @(*) begin
    DBusCachedPlugin_exceptionBus_valid = 1'b0;
    if(when_DBusCachedPlugin_l446) begin
      if(dataCache_1_io_cpu_writeBack_accessError) begin
        DBusCachedPlugin_exceptionBus_valid = 1'b1;
      end
      if(dataCache_1_io_cpu_writeBack_mmuException) begin
        DBusCachedPlugin_exceptionBus_valid = 1'b1;
      end
      if(dataCache_1_io_cpu_writeBack_unalignedAccess) begin
        DBusCachedPlugin_exceptionBus_valid = 1'b1;
      end
      if(dataCache_1_io_cpu_redo) begin
        DBusCachedPlugin_exceptionBus_valid = 1'b0;
      end
    end
  end

  assign DBusCachedPlugin_exceptionBus_payload_badAddr = writeBack_REGFILE_WRITE_DATA;
  always @(*) begin
    DBusCachedPlugin_exceptionBus_payload_code = 4'bxxxx;
    if(when_DBusCachedPlugin_l446) begin
      if(dataCache_1_io_cpu_writeBack_accessError) begin
        DBusCachedPlugin_exceptionBus_payload_code = {1'd0, _zz_DBusCachedPlugin_exceptionBus_payload_code};
      end
      if(dataCache_1_io_cpu_writeBack_mmuException) begin
        DBusCachedPlugin_exceptionBus_payload_code = (writeBack_MEMORY_WR ? 4'b1111 : 4'b1101);
      end
      if(dataCache_1_io_cpu_writeBack_unalignedAccess) begin
        DBusCachedPlugin_exceptionBus_payload_code = {1'd0, _zz_DBusCachedPlugin_exceptionBus_payload_code_1};
      end
    end
  end

  assign when_DBusCachedPlugin_l446 = (writeBack_arbitration_isValid && writeBack_MEMORY_ENABLE);
  assign when_DBusCachedPlugin_l466 = (dataCache_1_io_cpu_writeBack_isValid && dataCache_1_io_cpu_writeBack_haltIt);
  assign writeBack_DBusCachedPlugin_rspSplits_0 = dataCache_1_io_cpu_writeBack_data[7 : 0];
  assign writeBack_DBusCachedPlugin_rspSplits_1 = dataCache_1_io_cpu_writeBack_data[15 : 8];
  assign writeBack_DBusCachedPlugin_rspSplits_2 = dataCache_1_io_cpu_writeBack_data[23 : 16];
  assign writeBack_DBusCachedPlugin_rspSplits_3 = dataCache_1_io_cpu_writeBack_data[31 : 24];
  always @(*) begin
    writeBack_DBusCachedPlugin_rspShifted[7 : 0] = _zz_writeBack_DBusCachedPlugin_rspShifted;
    writeBack_DBusCachedPlugin_rspShifted[15 : 8] = _zz_writeBack_DBusCachedPlugin_rspShifted_2;
    writeBack_DBusCachedPlugin_rspShifted[23 : 16] = writeBack_DBusCachedPlugin_rspSplits_2;
    writeBack_DBusCachedPlugin_rspShifted[31 : 24] = writeBack_DBusCachedPlugin_rspSplits_3;
  end

  assign writeBack_DBusCachedPlugin_rspRf = writeBack_DBusCachedPlugin_rspShifted[31 : 0];
  assign switch_Misc_l210 = writeBack_INSTRUCTION[13 : 12];
  assign _zz_writeBack_DBusCachedPlugin_rspFormated = (writeBack_DBusCachedPlugin_rspRf[7] && (! writeBack_INSTRUCTION[14]));
  always @(*) begin
    _zz_writeBack_DBusCachedPlugin_rspFormated_1[31] = _zz_writeBack_DBusCachedPlugin_rspFormated;
    _zz_writeBack_DBusCachedPlugin_rspFormated_1[30] = _zz_writeBack_DBusCachedPlugin_rspFormated;
    _zz_writeBack_DBusCachedPlugin_rspFormated_1[29] = _zz_writeBack_DBusCachedPlugin_rspFormated;
    _zz_writeBack_DBusCachedPlugin_rspFormated_1[28] = _zz_writeBack_DBusCachedPlugin_rspFormated;
    _zz_writeBack_DBusCachedPlugin_rspFormated_1[27] = _zz_writeBack_DBusCachedPlugin_rspFormated;
    _zz_writeBack_DBusCachedPlugin_rspFormated_1[26] = _zz_writeBack_DBusCachedPlugin_rspFormated;
    _zz_writeBack_DBusCachedPlugin_rspFormated_1[25] = _zz_writeBack_DBusCachedPlugin_rspFormated;
    _zz_writeBack_DBusCachedPlugin_rspFormated_1[24] = _zz_writeBack_DBusCachedPlugin_rspFormated;
    _zz_writeBack_DBusCachedPlugin_rspFormated_1[23] = _zz_writeBack_DBusCachedPlugin_rspFormated;
    _zz_writeBack_DBusCachedPlugin_rspFormated_1[22] = _zz_writeBack_DBusCachedPlugin_rspFormated;
    _zz_writeBack_DBusCachedPlugin_rspFormated_1[21] = _zz_writeBack_DBusCachedPlugin_rspFormated;
    _zz_writeBack_DBusCachedPlugin_rspFormated_1[20] = _zz_writeBack_DBusCachedPlugin_rspFormated;
    _zz_writeBack_DBusCachedPlugin_rspFormated_1[19] = _zz_writeBack_DBusCachedPlugin_rspFormated;
    _zz_writeBack_DBusCachedPlugin_rspFormated_1[18] = _zz_writeBack_DBusCachedPlugin_rspFormated;
    _zz_writeBack_DBusCachedPlugin_rspFormated_1[17] = _zz_writeBack_DBusCachedPlugin_rspFormated;
    _zz_writeBack_DBusCachedPlugin_rspFormated_1[16] = _zz_writeBack_DBusCachedPlugin_rspFormated;
    _zz_writeBack_DBusCachedPlugin_rspFormated_1[15] = _zz_writeBack_DBusCachedPlugin_rspFormated;
    _zz_writeBack_DBusCachedPlugin_rspFormated_1[14] = _zz_writeBack_DBusCachedPlugin_rspFormated;
    _zz_writeBack_DBusCachedPlugin_rspFormated_1[13] = _zz_writeBack_DBusCachedPlugin_rspFormated;
    _zz_writeBack_DBusCachedPlugin_rspFormated_1[12] = _zz_writeBack_DBusCachedPlugin_rspFormated;
    _zz_writeBack_DBusCachedPlugin_rspFormated_1[11] = _zz_writeBack_DBusCachedPlugin_rspFormated;
    _zz_writeBack_DBusCachedPlugin_rspFormated_1[10] = _zz_writeBack_DBusCachedPlugin_rspFormated;
    _zz_writeBack_DBusCachedPlugin_rspFormated_1[9] = _zz_writeBack_DBusCachedPlugin_rspFormated;
    _zz_writeBack_DBusCachedPlugin_rspFormated_1[8] = _zz_writeBack_DBusCachedPlugin_rspFormated;
    _zz_writeBack_DBusCachedPlugin_rspFormated_1[7 : 0] = writeBack_DBusCachedPlugin_rspRf[7 : 0];
  end

  assign _zz_writeBack_DBusCachedPlugin_rspFormated_2 = (writeBack_DBusCachedPlugin_rspRf[15] && (! writeBack_INSTRUCTION[14]));
  always @(*) begin
    _zz_writeBack_DBusCachedPlugin_rspFormated_3[31] = _zz_writeBack_DBusCachedPlugin_rspFormated_2;
    _zz_writeBack_DBusCachedPlugin_rspFormated_3[30] = _zz_writeBack_DBusCachedPlugin_rspFormated_2;
    _zz_writeBack_DBusCachedPlugin_rspFormated_3[29] = _zz_writeBack_DBusCachedPlugin_rspFormated_2;
    _zz_writeBack_DBusCachedPlugin_rspFormated_3[28] = _zz_writeBack_DBusCachedPlugin_rspFormated_2;
    _zz_writeBack_DBusCachedPlugin_rspFormated_3[27] = _zz_writeBack_DBusCachedPlugin_rspFormated_2;
    _zz_writeBack_DBusCachedPlugin_rspFormated_3[26] = _zz_writeBack_DBusCachedPlugin_rspFormated_2;
    _zz_writeBack_DBusCachedPlugin_rspFormated_3[25] = _zz_writeBack_DBusCachedPlugin_rspFormated_2;
    _zz_writeBack_DBusCachedPlugin_rspFormated_3[24] = _zz_writeBack_DBusCachedPlugin_rspFormated_2;
    _zz_writeBack_DBusCachedPlugin_rspFormated_3[23] = _zz_writeBack_DBusCachedPlugin_rspFormated_2;
    _zz_writeBack_DBusCachedPlugin_rspFormated_3[22] = _zz_writeBack_DBusCachedPlugin_rspFormated_2;
    _zz_writeBack_DBusCachedPlugin_rspFormated_3[21] = _zz_writeBack_DBusCachedPlugin_rspFormated_2;
    _zz_writeBack_DBusCachedPlugin_rspFormated_3[20] = _zz_writeBack_DBusCachedPlugin_rspFormated_2;
    _zz_writeBack_DBusCachedPlugin_rspFormated_3[19] = _zz_writeBack_DBusCachedPlugin_rspFormated_2;
    _zz_writeBack_DBusCachedPlugin_rspFormated_3[18] = _zz_writeBack_DBusCachedPlugin_rspFormated_2;
    _zz_writeBack_DBusCachedPlugin_rspFormated_3[17] = _zz_writeBack_DBusCachedPlugin_rspFormated_2;
    _zz_writeBack_DBusCachedPlugin_rspFormated_3[16] = _zz_writeBack_DBusCachedPlugin_rspFormated_2;
    _zz_writeBack_DBusCachedPlugin_rspFormated_3[15 : 0] = writeBack_DBusCachedPlugin_rspRf[15 : 0];
  end

  always @(*) begin
    case(switch_Misc_l210)
      2'b00 : begin
        writeBack_DBusCachedPlugin_rspFormated = _zz_writeBack_DBusCachedPlugin_rspFormated_1;
      end
      2'b01 : begin
        writeBack_DBusCachedPlugin_rspFormated = _zz_writeBack_DBusCachedPlugin_rspFormated_3;
      end
      default : begin
        writeBack_DBusCachedPlugin_rspFormated = writeBack_DBusCachedPlugin_rspRf;
      end
    endcase
  end

  assign when_DBusCachedPlugin_l492 = (writeBack_arbitration_isValid && writeBack_MEMORY_ENABLE);
  assign when_PmpPlugin_l138 = (! execute_arbitration_isStuck);
  always @(*) begin
    execute_PmpPlugin_fsmComplete = 1'b0;
    if(when_StateMachine_l249) begin
      execute_PmpPlugin_fsmComplete = 1'b1;
    end
  end

  assign execute_PmpPlugin_csrAddress = execute_INSTRUCTION[31 : 20];
  assign execute_PmpPlugin_pmpNcfg = execute_PmpPlugin_csrAddress[3 : 0];
  assign execute_PmpPlugin_pmpcfgN = execute_PmpPlugin_pmpNcfg[1 : 0];
  assign execute_PmpPlugin_pmpcfgCsr = (execute_INSTRUCTION[31 : 24] == 8'h3a);
  assign execute_PmpPlugin_pmpaddrCsr = (execute_INSTRUCTION[31 : 24] == 8'h3b);
  assign execute_PmpPlugin_fsm_wantExit = 1'b0;
  always @(*) begin
    execute_PmpPlugin_fsm_wantStart = 1'b0;
    case(execute_PmpPlugin_fsm_stateReg)
      execute_PmpPlugin_fsm_enumDef_stateIdle : begin
      end
      execute_PmpPlugin_fsm_enumDef_stateWrite : begin
      end
      execute_PmpPlugin_fsm_enumDef_stateCfg : begin
      end
      execute_PmpPlugin_fsm_enumDef_stateAddr : begin
      end
      default : begin
        execute_PmpPlugin_fsm_wantStart = 1'b1;
      end
    endcase
  end

  assign execute_PmpPlugin_fsm_wantKill = 1'b0;
  always @(*) begin
    if(execute_PmpPlugin_pmpaddrCsr_) begin
      PmpPlugin_setter_io_addr = execute_PmpPlugin_writeData_;
    end else begin
      PmpPlugin_setter_io_addr = _zz_PmpPlugin_pmpaddr_port0;
    end
  end

  assign when_PmpPlugin_l246 = (execute_PmpPlugin_fsm_fsmEnable && (! _zz_when_PmpPlugin_l246[7]));
  assign _zz_8 = ({15'd0,1'b1} <<< execute_PmpPlugin_fsm_fsmCounter);
  assign _zz_9 = ({15'd0,1'b1} <<< execute_PmpPlugin_fsm_fsmCounter);
  assign DBusCachedPlugin_mmuBus_rsp_physicalAddress = DBusCachedPlugin_mmuBus_cmd_0_virtualAddress;
  assign DBusCachedPlugin_mmuBus_rsp_isIoAccess = DBusCachedPlugin_mmuBus_cmd_0_virtualAddress[31];
  assign DBusCachedPlugin_mmuBus_rsp_isPaging = 1'b0;
  assign DBusCachedPlugin_mmuBus_rsp_exception = 1'b0;
  assign DBusCachedPlugin_mmuBus_rsp_refilling = 1'b0;
  assign DBusCachedPlugin_mmuBus_rsp_allowExecute = 1'b0;
  assign DBusCachedPlugin_mmuBus_busy = 1'b0;
  assign _zz_PmpPlugin_dGuard_hits_0 = DBusCachedPlugin_mmuBus_cmd_0_virtualAddress[31 : 7];
  assign PmpPlugin_dGuard_hits_0 = ((((_zz_PmpPlugin_dGuard_hits_0 & _zz_PmpPlugin_dGuard_hits_0_1) == _zz_PmpPlugin_dGuard_hits_0_3) && (PmpPlugin_pmpcfg_0[7] || (! (CsrPlugin_privilege == 2'b11)))) && (PmpPlugin_pmpcfg_0[4 : 3] == 2'b11));
  assign PmpPlugin_dGuard_hits_1 = ((((_zz_PmpPlugin_dGuard_hits_0 & _zz_PmpPlugin_dGuard_hits_1) == _zz_PmpPlugin_dGuard_hits_1_2) && (PmpPlugin_pmpcfg_1[7] || (! (CsrPlugin_privilege == 2'b11)))) && (PmpPlugin_pmpcfg_1[4 : 3] == 2'b11));
  assign PmpPlugin_dGuard_hits_2 = ((((_zz_PmpPlugin_dGuard_hits_0 & _zz_PmpPlugin_dGuard_hits_2) == _zz_PmpPlugin_dGuard_hits_2_2) && (PmpPlugin_pmpcfg_2[7] || (! (CsrPlugin_privilege == 2'b11)))) && (PmpPlugin_pmpcfg_2[4 : 3] == 2'b11));
  assign PmpPlugin_dGuard_hits_3 = ((((_zz_PmpPlugin_dGuard_hits_0 & _zz_PmpPlugin_dGuard_hits_3) == _zz_PmpPlugin_dGuard_hits_3_2) && (PmpPlugin_pmpcfg_3[7] || (! (CsrPlugin_privilege == 2'b11)))) && (PmpPlugin_pmpcfg_3[4 : 3] == 2'b11));
  assign PmpPlugin_dGuard_hits_4 = ((((_zz_PmpPlugin_dGuard_hits_0 & _zz_PmpPlugin_dGuard_hits_4) == _zz_PmpPlugin_dGuard_hits_4_2) && (PmpPlugin_pmpcfg_4[7] || (! (CsrPlugin_privilege == 2'b11)))) && (PmpPlugin_pmpcfg_4[4 : 3] == 2'b11));
  assign PmpPlugin_dGuard_hits_5 = ((((_zz_PmpPlugin_dGuard_hits_0 & _zz_PmpPlugin_dGuard_hits_5) == _zz_PmpPlugin_dGuard_hits_5_2) && (PmpPlugin_pmpcfg_5[7] || (! (CsrPlugin_privilege == 2'b11)))) && (PmpPlugin_pmpcfg_5[4 : 3] == 2'b11));
  assign PmpPlugin_dGuard_hits_6 = ((((_zz_PmpPlugin_dGuard_hits_0 & _zz_PmpPlugin_dGuard_hits_6) == _zz_PmpPlugin_dGuard_hits_6_2) && (PmpPlugin_pmpcfg_6[7] || (! (CsrPlugin_privilege == 2'b11)))) && (PmpPlugin_pmpcfg_6[4 : 3] == 2'b11));
  assign PmpPlugin_dGuard_hits_7 = ((((_zz_PmpPlugin_dGuard_hits_0 & _zz_PmpPlugin_dGuard_hits_7) == _zz_PmpPlugin_dGuard_hits_7_2) && (PmpPlugin_pmpcfg_7[7] || (! (CsrPlugin_privilege == 2'b11)))) && (PmpPlugin_pmpcfg_7[4 : 3] == 2'b11));
  assign PmpPlugin_dGuard_hits_8 = ((((_zz_PmpPlugin_dGuard_hits_0 & _zz_PmpPlugin_dGuard_hits_8) == _zz_PmpPlugin_dGuard_hits_8_2) && (PmpPlugin_pmpcfg_8[7] || (! (CsrPlugin_privilege == 2'b11)))) && (PmpPlugin_pmpcfg_8[4 : 3] == 2'b11));
  assign PmpPlugin_dGuard_hits_9 = ((((_zz_PmpPlugin_dGuard_hits_0 & _zz_PmpPlugin_dGuard_hits_9) == _zz_PmpPlugin_dGuard_hits_9_2) && (PmpPlugin_pmpcfg_9[7] || (! (CsrPlugin_privilege == 2'b11)))) && (PmpPlugin_pmpcfg_9[4 : 3] == 2'b11));
  assign PmpPlugin_dGuard_hits_10 = ((((_zz_PmpPlugin_dGuard_hits_0 & _zz_PmpPlugin_dGuard_hits_10) == _zz_PmpPlugin_dGuard_hits_10_2) && (PmpPlugin_pmpcfg_10[7] || (! (CsrPlugin_privilege == 2'b11)))) && (PmpPlugin_pmpcfg_10[4 : 3] == 2'b11));
  assign PmpPlugin_dGuard_hits_11 = ((((_zz_PmpPlugin_dGuard_hits_0 & _zz_PmpPlugin_dGuard_hits_11) == _zz_PmpPlugin_dGuard_hits_11_2) && (PmpPlugin_pmpcfg_11[7] || (! (CsrPlugin_privilege == 2'b11)))) && (PmpPlugin_pmpcfg_11[4 : 3] == 2'b11));
  assign PmpPlugin_dGuard_hits_12 = ((((_zz_PmpPlugin_dGuard_hits_0 & _zz_PmpPlugin_dGuard_hits_12) == _zz_PmpPlugin_dGuard_hits_12_2) && (PmpPlugin_pmpcfg_12[7] || (! (CsrPlugin_privilege == 2'b11)))) && (PmpPlugin_pmpcfg_12[4 : 3] == 2'b11));
  assign PmpPlugin_dGuard_hits_13 = ((((_zz_PmpPlugin_dGuard_hits_0 & _zz_PmpPlugin_dGuard_hits_13) == _zz_PmpPlugin_dGuard_hits_13_2) && (PmpPlugin_pmpcfg_13[7] || (! (CsrPlugin_privilege == 2'b11)))) && (PmpPlugin_pmpcfg_13[4 : 3] == 2'b11));
  assign PmpPlugin_dGuard_hits_14 = ((((_zz_PmpPlugin_dGuard_hits_0 & _zz_PmpPlugin_dGuard_hits_14) == _zz_PmpPlugin_dGuard_hits_14_2) && (PmpPlugin_pmpcfg_14[7] || (! (CsrPlugin_privilege == 2'b11)))) && (PmpPlugin_pmpcfg_14[4 : 3] == 2'b11));
  assign PmpPlugin_dGuard_hits_15 = ((((_zz_PmpPlugin_dGuard_hits_0 & _zz_PmpPlugin_dGuard_hits_15) == _zz_PmpPlugin_dGuard_hits_15_2) && (PmpPlugin_pmpcfg_15[7] || (! (CsrPlugin_privilege == 2'b11)))) && (PmpPlugin_pmpcfg_15[4 : 3] == 2'b11));
  assign when_PmpPlugin_l277 = (! ({PmpPlugin_dGuard_hits_15,{PmpPlugin_dGuard_hits_14,{PmpPlugin_dGuard_hits_13,{PmpPlugin_dGuard_hits_12,{PmpPlugin_dGuard_hits_11,{PmpPlugin_dGuard_hits_10,{PmpPlugin_dGuard_hits_9,{PmpPlugin_dGuard_hits_8,{PmpPlugin_dGuard_hits_7,{_zz_when_PmpPlugin_l277,_zz_when_PmpPlugin_l277_1}}}}}}}}}} != 16'h0));
  always @(*) begin
    if(when_PmpPlugin_l277) begin
      DBusCachedPlugin_mmuBus_rsp_allowRead = (CsrPlugin_privilege == 2'b11);
    end else begin
      DBusCachedPlugin_mmuBus_rsp_allowRead = _zz_DBusCachedPlugin_mmuBus_rsp_allowRead_17;
    end
  end

  always @(*) begin
    if(when_PmpPlugin_l277) begin
      DBusCachedPlugin_mmuBus_rsp_allowWrite = (CsrPlugin_privilege == 2'b11);
    end else begin
      DBusCachedPlugin_mmuBus_rsp_allowWrite = _zz_DBusCachedPlugin_mmuBus_rsp_allowWrite_17;
    end
  end

  assign _zz_DBusCachedPlugin_mmuBus_rsp_allowRead = {PmpPlugin_dGuard_hits_15,{PmpPlugin_dGuard_hits_14,{PmpPlugin_dGuard_hits_13,{PmpPlugin_dGuard_hits_12,{PmpPlugin_dGuard_hits_11,{PmpPlugin_dGuard_hits_10,{PmpPlugin_dGuard_hits_9,{PmpPlugin_dGuard_hits_8,{PmpPlugin_dGuard_hits_7,{PmpPlugin_dGuard_hits_6,{_zz__zz_DBusCachedPlugin_mmuBus_rsp_allowRead,_zz__zz_DBusCachedPlugin_mmuBus_rsp_allowRead_1}}}}}}}}}}};
  assign _zz_DBusCachedPlugin_mmuBus_rsp_allowRead_1 = (_zz_DBusCachedPlugin_mmuBus_rsp_allowRead & (~ _zz__zz_DBusCachedPlugin_mmuBus_rsp_allowRead_1_1));
  assign _zz_DBusCachedPlugin_mmuBus_rsp_allowRead_2 = _zz_DBusCachedPlugin_mmuBus_rsp_allowRead_1[3];
  assign _zz_DBusCachedPlugin_mmuBus_rsp_allowRead_3 = _zz_DBusCachedPlugin_mmuBus_rsp_allowRead_1[5];
  assign _zz_DBusCachedPlugin_mmuBus_rsp_allowRead_4 = _zz_DBusCachedPlugin_mmuBus_rsp_allowRead_1[6];
  assign _zz_DBusCachedPlugin_mmuBus_rsp_allowRead_5 = _zz_DBusCachedPlugin_mmuBus_rsp_allowRead_1[7];
  assign _zz_DBusCachedPlugin_mmuBus_rsp_allowRead_6 = _zz_DBusCachedPlugin_mmuBus_rsp_allowRead_1[9];
  assign _zz_DBusCachedPlugin_mmuBus_rsp_allowRead_7 = _zz_DBusCachedPlugin_mmuBus_rsp_allowRead_1[10];
  assign _zz_DBusCachedPlugin_mmuBus_rsp_allowRead_8 = _zz_DBusCachedPlugin_mmuBus_rsp_allowRead_1[11];
  assign _zz_DBusCachedPlugin_mmuBus_rsp_allowRead_9 = _zz_DBusCachedPlugin_mmuBus_rsp_allowRead_1[12];
  assign _zz_DBusCachedPlugin_mmuBus_rsp_allowRead_10 = _zz_DBusCachedPlugin_mmuBus_rsp_allowRead_1[13];
  assign _zz_DBusCachedPlugin_mmuBus_rsp_allowRead_11 = _zz_DBusCachedPlugin_mmuBus_rsp_allowRead_1[14];
  assign _zz_DBusCachedPlugin_mmuBus_rsp_allowRead_12 = _zz_DBusCachedPlugin_mmuBus_rsp_allowRead_1[15];
  assign _zz_DBusCachedPlugin_mmuBus_rsp_allowRead_13 = (((((((_zz_DBusCachedPlugin_mmuBus_rsp_allowRead_1[1] || _zz_DBusCachedPlugin_mmuBus_rsp_allowRead_2) || _zz_DBusCachedPlugin_mmuBus_rsp_allowRead_3) || _zz_DBusCachedPlugin_mmuBus_rsp_allowRead_5) || _zz_DBusCachedPlugin_mmuBus_rsp_allowRead_6) || _zz_DBusCachedPlugin_mmuBus_rsp_allowRead_8) || _zz_DBusCachedPlugin_mmuBus_rsp_allowRead_10) || _zz_DBusCachedPlugin_mmuBus_rsp_allowRead_12);
  assign _zz_DBusCachedPlugin_mmuBus_rsp_allowRead_14 = (((((((_zz_DBusCachedPlugin_mmuBus_rsp_allowRead_1[2] || _zz_DBusCachedPlugin_mmuBus_rsp_allowRead_2) || _zz_DBusCachedPlugin_mmuBus_rsp_allowRead_4) || _zz_DBusCachedPlugin_mmuBus_rsp_allowRead_5) || _zz_DBusCachedPlugin_mmuBus_rsp_allowRead_7) || _zz_DBusCachedPlugin_mmuBus_rsp_allowRead_8) || _zz_DBusCachedPlugin_mmuBus_rsp_allowRead_11) || _zz_DBusCachedPlugin_mmuBus_rsp_allowRead_12);
  assign _zz_DBusCachedPlugin_mmuBus_rsp_allowRead_15 = (((((((_zz_DBusCachedPlugin_mmuBus_rsp_allowRead_1[4] || _zz_DBusCachedPlugin_mmuBus_rsp_allowRead_3) || _zz_DBusCachedPlugin_mmuBus_rsp_allowRead_4) || _zz_DBusCachedPlugin_mmuBus_rsp_allowRead_5) || _zz_DBusCachedPlugin_mmuBus_rsp_allowRead_9) || _zz_DBusCachedPlugin_mmuBus_rsp_allowRead_10) || _zz_DBusCachedPlugin_mmuBus_rsp_allowRead_11) || _zz_DBusCachedPlugin_mmuBus_rsp_allowRead_12);
  assign _zz_DBusCachedPlugin_mmuBus_rsp_allowRead_16 = (((((((_zz_DBusCachedPlugin_mmuBus_rsp_allowRead_1[8] || _zz_DBusCachedPlugin_mmuBus_rsp_allowRead_6) || _zz_DBusCachedPlugin_mmuBus_rsp_allowRead_7) || _zz_DBusCachedPlugin_mmuBus_rsp_allowRead_8) || _zz_DBusCachedPlugin_mmuBus_rsp_allowRead_9) || _zz_DBusCachedPlugin_mmuBus_rsp_allowRead_10) || _zz_DBusCachedPlugin_mmuBus_rsp_allowRead_11) || _zz_DBusCachedPlugin_mmuBus_rsp_allowRead_12);
  assign _zz_DBusCachedPlugin_mmuBus_rsp_allowWrite = {PmpPlugin_dGuard_hits_15,{PmpPlugin_dGuard_hits_14,{PmpPlugin_dGuard_hits_13,{PmpPlugin_dGuard_hits_12,{PmpPlugin_dGuard_hits_11,{PmpPlugin_dGuard_hits_10,{PmpPlugin_dGuard_hits_9,{PmpPlugin_dGuard_hits_8,{PmpPlugin_dGuard_hits_7,{PmpPlugin_dGuard_hits_6,{_zz__zz_DBusCachedPlugin_mmuBus_rsp_allowWrite,_zz__zz_DBusCachedPlugin_mmuBus_rsp_allowWrite_1}}}}}}}}}}};
  assign _zz_DBusCachedPlugin_mmuBus_rsp_allowWrite_1 = (_zz_DBusCachedPlugin_mmuBus_rsp_allowWrite & (~ _zz__zz_DBusCachedPlugin_mmuBus_rsp_allowWrite_1_1));
  assign _zz_DBusCachedPlugin_mmuBus_rsp_allowWrite_2 = _zz_DBusCachedPlugin_mmuBus_rsp_allowWrite_1[3];
  assign _zz_DBusCachedPlugin_mmuBus_rsp_allowWrite_3 = _zz_DBusCachedPlugin_mmuBus_rsp_allowWrite_1[5];
  assign _zz_DBusCachedPlugin_mmuBus_rsp_allowWrite_4 = _zz_DBusCachedPlugin_mmuBus_rsp_allowWrite_1[6];
  assign _zz_DBusCachedPlugin_mmuBus_rsp_allowWrite_5 = _zz_DBusCachedPlugin_mmuBus_rsp_allowWrite_1[7];
  assign _zz_DBusCachedPlugin_mmuBus_rsp_allowWrite_6 = _zz_DBusCachedPlugin_mmuBus_rsp_allowWrite_1[9];
  assign _zz_DBusCachedPlugin_mmuBus_rsp_allowWrite_7 = _zz_DBusCachedPlugin_mmuBus_rsp_allowWrite_1[10];
  assign _zz_DBusCachedPlugin_mmuBus_rsp_allowWrite_8 = _zz_DBusCachedPlugin_mmuBus_rsp_allowWrite_1[11];
  assign _zz_DBusCachedPlugin_mmuBus_rsp_allowWrite_9 = _zz_DBusCachedPlugin_mmuBus_rsp_allowWrite_1[12];
  assign _zz_DBusCachedPlugin_mmuBus_rsp_allowWrite_10 = _zz_DBusCachedPlugin_mmuBus_rsp_allowWrite_1[13];
  assign _zz_DBusCachedPlugin_mmuBus_rsp_allowWrite_11 = _zz_DBusCachedPlugin_mmuBus_rsp_allowWrite_1[14];
  assign _zz_DBusCachedPlugin_mmuBus_rsp_allowWrite_12 = _zz_DBusCachedPlugin_mmuBus_rsp_allowWrite_1[15];
  assign _zz_DBusCachedPlugin_mmuBus_rsp_allowWrite_13 = (((((((_zz_DBusCachedPlugin_mmuBus_rsp_allowWrite_1[1] || _zz_DBusCachedPlugin_mmuBus_rsp_allowWrite_2) || _zz_DBusCachedPlugin_mmuBus_rsp_allowWrite_3) || _zz_DBusCachedPlugin_mmuBus_rsp_allowWrite_5) || _zz_DBusCachedPlugin_mmuBus_rsp_allowWrite_6) || _zz_DBusCachedPlugin_mmuBus_rsp_allowWrite_8) || _zz_DBusCachedPlugin_mmuBus_rsp_allowWrite_10) || _zz_DBusCachedPlugin_mmuBus_rsp_allowWrite_12);
  assign _zz_DBusCachedPlugin_mmuBus_rsp_allowWrite_14 = (((((((_zz_DBusCachedPlugin_mmuBus_rsp_allowWrite_1[2] || _zz_DBusCachedPlugin_mmuBus_rsp_allowWrite_2) || _zz_DBusCachedPlugin_mmuBus_rsp_allowWrite_4) || _zz_DBusCachedPlugin_mmuBus_rsp_allowWrite_5) || _zz_DBusCachedPlugin_mmuBus_rsp_allowWrite_7) || _zz_DBusCachedPlugin_mmuBus_rsp_allowWrite_8) || _zz_DBusCachedPlugin_mmuBus_rsp_allowWrite_11) || _zz_DBusCachedPlugin_mmuBus_rsp_allowWrite_12);
  assign _zz_DBusCachedPlugin_mmuBus_rsp_allowWrite_15 = (((((((_zz_DBusCachedPlugin_mmuBus_rsp_allowWrite_1[4] || _zz_DBusCachedPlugin_mmuBus_rsp_allowWrite_3) || _zz_DBusCachedPlugin_mmuBus_rsp_allowWrite_4) || _zz_DBusCachedPlugin_mmuBus_rsp_allowWrite_5) || _zz_DBusCachedPlugin_mmuBus_rsp_allowWrite_9) || _zz_DBusCachedPlugin_mmuBus_rsp_allowWrite_10) || _zz_DBusCachedPlugin_mmuBus_rsp_allowWrite_11) || _zz_DBusCachedPlugin_mmuBus_rsp_allowWrite_12);
  assign _zz_DBusCachedPlugin_mmuBus_rsp_allowWrite_16 = (((((((_zz_DBusCachedPlugin_mmuBus_rsp_allowWrite_1[8] || _zz_DBusCachedPlugin_mmuBus_rsp_allowWrite_6) || _zz_DBusCachedPlugin_mmuBus_rsp_allowWrite_7) || _zz_DBusCachedPlugin_mmuBus_rsp_allowWrite_8) || _zz_DBusCachedPlugin_mmuBus_rsp_allowWrite_9) || _zz_DBusCachedPlugin_mmuBus_rsp_allowWrite_10) || _zz_DBusCachedPlugin_mmuBus_rsp_allowWrite_11) || _zz_DBusCachedPlugin_mmuBus_rsp_allowWrite_12);
  assign IBusCachedPlugin_mmuBus_rsp_physicalAddress = IBusCachedPlugin_mmuBus_cmd_0_virtualAddress;
  assign IBusCachedPlugin_mmuBus_rsp_isIoAccess = IBusCachedPlugin_mmuBus_cmd_0_virtualAddress[31];
  assign IBusCachedPlugin_mmuBus_rsp_isPaging = 1'b0;
  assign IBusCachedPlugin_mmuBus_rsp_exception = 1'b0;
  assign IBusCachedPlugin_mmuBus_rsp_refilling = 1'b0;
  assign IBusCachedPlugin_mmuBus_rsp_allowRead = 1'b0;
  assign IBusCachedPlugin_mmuBus_rsp_allowWrite = 1'b0;
  assign IBusCachedPlugin_mmuBus_busy = 1'b0;
  assign _zz_PmpPlugin_iGuard_hits_0 = IBusCachedPlugin_mmuBus_cmd_0_virtualAddress[31 : 7];
  assign PmpPlugin_iGuard_hits_0 = ((((_zz_PmpPlugin_iGuard_hits_0 & _zz_PmpPlugin_iGuard_hits_0_1) == _zz_PmpPlugin_iGuard_hits_0_3) && (PmpPlugin_pmpcfg_0[7] || (! (CsrPlugin_privilege == 2'b11)))) && (PmpPlugin_pmpcfg_0[4 : 3] == 2'b11));
  assign PmpPlugin_iGuard_hits_1 = ((((_zz_PmpPlugin_iGuard_hits_0 & _zz_PmpPlugin_iGuard_hits_1) == _zz_PmpPlugin_iGuard_hits_1_2) && (PmpPlugin_pmpcfg_1[7] || (! (CsrPlugin_privilege == 2'b11)))) && (PmpPlugin_pmpcfg_1[4 : 3] == 2'b11));
  assign PmpPlugin_iGuard_hits_2 = ((((_zz_PmpPlugin_iGuard_hits_0 & _zz_PmpPlugin_iGuard_hits_2) == _zz_PmpPlugin_iGuard_hits_2_2) && (PmpPlugin_pmpcfg_2[7] || (! (CsrPlugin_privilege == 2'b11)))) && (PmpPlugin_pmpcfg_2[4 : 3] == 2'b11));
  assign PmpPlugin_iGuard_hits_3 = ((((_zz_PmpPlugin_iGuard_hits_0 & _zz_PmpPlugin_iGuard_hits_3) == _zz_PmpPlugin_iGuard_hits_3_2) && (PmpPlugin_pmpcfg_3[7] || (! (CsrPlugin_privilege == 2'b11)))) && (PmpPlugin_pmpcfg_3[4 : 3] == 2'b11));
  assign PmpPlugin_iGuard_hits_4 = ((((_zz_PmpPlugin_iGuard_hits_0 & _zz_PmpPlugin_iGuard_hits_4) == _zz_PmpPlugin_iGuard_hits_4_2) && (PmpPlugin_pmpcfg_4[7] || (! (CsrPlugin_privilege == 2'b11)))) && (PmpPlugin_pmpcfg_4[4 : 3] == 2'b11));
  assign PmpPlugin_iGuard_hits_5 = ((((_zz_PmpPlugin_iGuard_hits_0 & _zz_PmpPlugin_iGuard_hits_5) == _zz_PmpPlugin_iGuard_hits_5_2) && (PmpPlugin_pmpcfg_5[7] || (! (CsrPlugin_privilege == 2'b11)))) && (PmpPlugin_pmpcfg_5[4 : 3] == 2'b11));
  assign PmpPlugin_iGuard_hits_6 = ((((_zz_PmpPlugin_iGuard_hits_0 & _zz_PmpPlugin_iGuard_hits_6) == _zz_PmpPlugin_iGuard_hits_6_2) && (PmpPlugin_pmpcfg_6[7] || (! (CsrPlugin_privilege == 2'b11)))) && (PmpPlugin_pmpcfg_6[4 : 3] == 2'b11));
  assign PmpPlugin_iGuard_hits_7 = ((((_zz_PmpPlugin_iGuard_hits_0 & _zz_PmpPlugin_iGuard_hits_7) == _zz_PmpPlugin_iGuard_hits_7_2) && (PmpPlugin_pmpcfg_7[7] || (! (CsrPlugin_privilege == 2'b11)))) && (PmpPlugin_pmpcfg_7[4 : 3] == 2'b11));
  assign PmpPlugin_iGuard_hits_8 = ((((_zz_PmpPlugin_iGuard_hits_0 & _zz_PmpPlugin_iGuard_hits_8) == _zz_PmpPlugin_iGuard_hits_8_2) && (PmpPlugin_pmpcfg_8[7] || (! (CsrPlugin_privilege == 2'b11)))) && (PmpPlugin_pmpcfg_8[4 : 3] == 2'b11));
  assign PmpPlugin_iGuard_hits_9 = ((((_zz_PmpPlugin_iGuard_hits_0 & _zz_PmpPlugin_iGuard_hits_9) == _zz_PmpPlugin_iGuard_hits_9_2) && (PmpPlugin_pmpcfg_9[7] || (! (CsrPlugin_privilege == 2'b11)))) && (PmpPlugin_pmpcfg_9[4 : 3] == 2'b11));
  assign PmpPlugin_iGuard_hits_10 = ((((_zz_PmpPlugin_iGuard_hits_0 & _zz_PmpPlugin_iGuard_hits_10) == _zz_PmpPlugin_iGuard_hits_10_2) && (PmpPlugin_pmpcfg_10[7] || (! (CsrPlugin_privilege == 2'b11)))) && (PmpPlugin_pmpcfg_10[4 : 3] == 2'b11));
  assign PmpPlugin_iGuard_hits_11 = ((((_zz_PmpPlugin_iGuard_hits_0 & _zz_PmpPlugin_iGuard_hits_11) == _zz_PmpPlugin_iGuard_hits_11_2) && (PmpPlugin_pmpcfg_11[7] || (! (CsrPlugin_privilege == 2'b11)))) && (PmpPlugin_pmpcfg_11[4 : 3] == 2'b11));
  assign PmpPlugin_iGuard_hits_12 = ((((_zz_PmpPlugin_iGuard_hits_0 & _zz_PmpPlugin_iGuard_hits_12) == _zz_PmpPlugin_iGuard_hits_12_2) && (PmpPlugin_pmpcfg_12[7] || (! (CsrPlugin_privilege == 2'b11)))) && (PmpPlugin_pmpcfg_12[4 : 3] == 2'b11));
  assign PmpPlugin_iGuard_hits_13 = ((((_zz_PmpPlugin_iGuard_hits_0 & _zz_PmpPlugin_iGuard_hits_13) == _zz_PmpPlugin_iGuard_hits_13_2) && (PmpPlugin_pmpcfg_13[7] || (! (CsrPlugin_privilege == 2'b11)))) && (PmpPlugin_pmpcfg_13[4 : 3] == 2'b11));
  assign PmpPlugin_iGuard_hits_14 = ((((_zz_PmpPlugin_iGuard_hits_0 & _zz_PmpPlugin_iGuard_hits_14) == _zz_PmpPlugin_iGuard_hits_14_2) && (PmpPlugin_pmpcfg_14[7] || (! (CsrPlugin_privilege == 2'b11)))) && (PmpPlugin_pmpcfg_14[4 : 3] == 2'b11));
  assign PmpPlugin_iGuard_hits_15 = ((((_zz_PmpPlugin_iGuard_hits_0 & _zz_PmpPlugin_iGuard_hits_15) == _zz_PmpPlugin_iGuard_hits_15_2) && (PmpPlugin_pmpcfg_15[7] || (! (CsrPlugin_privilege == 2'b11)))) && (PmpPlugin_pmpcfg_15[4 : 3] == 2'b11));
  assign when_PmpPlugin_l299 = (! ({PmpPlugin_iGuard_hits_15,{PmpPlugin_iGuard_hits_14,{PmpPlugin_iGuard_hits_13,{PmpPlugin_iGuard_hits_12,{PmpPlugin_iGuard_hits_11,{PmpPlugin_iGuard_hits_10,{PmpPlugin_iGuard_hits_9,{PmpPlugin_iGuard_hits_8,{PmpPlugin_iGuard_hits_7,{_zz_when_PmpPlugin_l299,_zz_when_PmpPlugin_l299_1}}}}}}}}}} != 16'h0));
  always @(*) begin
    if(when_PmpPlugin_l299) begin
      IBusCachedPlugin_mmuBus_rsp_allowExecute = (CsrPlugin_privilege == 2'b11);
    end else begin
      IBusCachedPlugin_mmuBus_rsp_allowExecute = _zz_IBusCachedPlugin_mmuBus_rsp_allowExecute_17;
    end
  end

  assign _zz_IBusCachedPlugin_mmuBus_rsp_allowExecute = {PmpPlugin_iGuard_hits_15,{PmpPlugin_iGuard_hits_14,{PmpPlugin_iGuard_hits_13,{PmpPlugin_iGuard_hits_12,{PmpPlugin_iGuard_hits_11,{PmpPlugin_iGuard_hits_10,{PmpPlugin_iGuard_hits_9,{PmpPlugin_iGuard_hits_8,{PmpPlugin_iGuard_hits_7,{PmpPlugin_iGuard_hits_6,{_zz__zz_IBusCachedPlugin_mmuBus_rsp_allowExecute,_zz__zz_IBusCachedPlugin_mmuBus_rsp_allowExecute_1}}}}}}}}}}};
  assign _zz_IBusCachedPlugin_mmuBus_rsp_allowExecute_1 = (_zz_IBusCachedPlugin_mmuBus_rsp_allowExecute & (~ _zz__zz_IBusCachedPlugin_mmuBus_rsp_allowExecute_1_1));
  assign _zz_IBusCachedPlugin_mmuBus_rsp_allowExecute_2 = _zz_IBusCachedPlugin_mmuBus_rsp_allowExecute_1[3];
  assign _zz_IBusCachedPlugin_mmuBus_rsp_allowExecute_3 = _zz_IBusCachedPlugin_mmuBus_rsp_allowExecute_1[5];
  assign _zz_IBusCachedPlugin_mmuBus_rsp_allowExecute_4 = _zz_IBusCachedPlugin_mmuBus_rsp_allowExecute_1[6];
  assign _zz_IBusCachedPlugin_mmuBus_rsp_allowExecute_5 = _zz_IBusCachedPlugin_mmuBus_rsp_allowExecute_1[7];
  assign _zz_IBusCachedPlugin_mmuBus_rsp_allowExecute_6 = _zz_IBusCachedPlugin_mmuBus_rsp_allowExecute_1[9];
  assign _zz_IBusCachedPlugin_mmuBus_rsp_allowExecute_7 = _zz_IBusCachedPlugin_mmuBus_rsp_allowExecute_1[10];
  assign _zz_IBusCachedPlugin_mmuBus_rsp_allowExecute_8 = _zz_IBusCachedPlugin_mmuBus_rsp_allowExecute_1[11];
  assign _zz_IBusCachedPlugin_mmuBus_rsp_allowExecute_9 = _zz_IBusCachedPlugin_mmuBus_rsp_allowExecute_1[12];
  assign _zz_IBusCachedPlugin_mmuBus_rsp_allowExecute_10 = _zz_IBusCachedPlugin_mmuBus_rsp_allowExecute_1[13];
  assign _zz_IBusCachedPlugin_mmuBus_rsp_allowExecute_11 = _zz_IBusCachedPlugin_mmuBus_rsp_allowExecute_1[14];
  assign _zz_IBusCachedPlugin_mmuBus_rsp_allowExecute_12 = _zz_IBusCachedPlugin_mmuBus_rsp_allowExecute_1[15];
  assign _zz_IBusCachedPlugin_mmuBus_rsp_allowExecute_13 = (((((((_zz_IBusCachedPlugin_mmuBus_rsp_allowExecute_1[1] || _zz_IBusCachedPlugin_mmuBus_rsp_allowExecute_2) || _zz_IBusCachedPlugin_mmuBus_rsp_allowExecute_3) || _zz_IBusCachedPlugin_mmuBus_rsp_allowExecute_5) || _zz_IBusCachedPlugin_mmuBus_rsp_allowExecute_6) || _zz_IBusCachedPlugin_mmuBus_rsp_allowExecute_8) || _zz_IBusCachedPlugin_mmuBus_rsp_allowExecute_10) || _zz_IBusCachedPlugin_mmuBus_rsp_allowExecute_12);
  assign _zz_IBusCachedPlugin_mmuBus_rsp_allowExecute_14 = (((((((_zz_IBusCachedPlugin_mmuBus_rsp_allowExecute_1[2] || _zz_IBusCachedPlugin_mmuBus_rsp_allowExecute_2) || _zz_IBusCachedPlugin_mmuBus_rsp_allowExecute_4) || _zz_IBusCachedPlugin_mmuBus_rsp_allowExecute_5) || _zz_IBusCachedPlugin_mmuBus_rsp_allowExecute_7) || _zz_IBusCachedPlugin_mmuBus_rsp_allowExecute_8) || _zz_IBusCachedPlugin_mmuBus_rsp_allowExecute_11) || _zz_IBusCachedPlugin_mmuBus_rsp_allowExecute_12);
  assign _zz_IBusCachedPlugin_mmuBus_rsp_allowExecute_15 = (((((((_zz_IBusCachedPlugin_mmuBus_rsp_allowExecute_1[4] || _zz_IBusCachedPlugin_mmuBus_rsp_allowExecute_3) || _zz_IBusCachedPlugin_mmuBus_rsp_allowExecute_4) || _zz_IBusCachedPlugin_mmuBus_rsp_allowExecute_5) || _zz_IBusCachedPlugin_mmuBus_rsp_allowExecute_9) || _zz_IBusCachedPlugin_mmuBus_rsp_allowExecute_10) || _zz_IBusCachedPlugin_mmuBus_rsp_allowExecute_11) || _zz_IBusCachedPlugin_mmuBus_rsp_allowExecute_12);
  assign _zz_IBusCachedPlugin_mmuBus_rsp_allowExecute_16 = (((((((_zz_IBusCachedPlugin_mmuBus_rsp_allowExecute_1[8] || _zz_IBusCachedPlugin_mmuBus_rsp_allowExecute_6) || _zz_IBusCachedPlugin_mmuBus_rsp_allowExecute_7) || _zz_IBusCachedPlugin_mmuBus_rsp_allowExecute_8) || _zz_IBusCachedPlugin_mmuBus_rsp_allowExecute_9) || _zz_IBusCachedPlugin_mmuBus_rsp_allowExecute_10) || _zz_IBusCachedPlugin_mmuBus_rsp_allowExecute_11) || _zz_IBusCachedPlugin_mmuBus_rsp_allowExecute_12);
  assign _zz_decode_IS_RS2_SIGNED_1 = ((decode_INSTRUCTION & 32'h00004050) == 32'h00004050);
  assign _zz_decode_IS_RS2_SIGNED_2 = ((decode_INSTRUCTION & 32'h00000018) == 32'h0);
  assign _zz_decode_IS_RS2_SIGNED_3 = ((decode_INSTRUCTION & 32'h00000004) == 32'h00000004);
  assign _zz_decode_IS_RS2_SIGNED_4 = ((decode_INSTRUCTION & 32'h00000048) == 32'h00000048);
  assign _zz_decode_IS_RS2_SIGNED_5 = ((decode_INSTRUCTION & 32'h00001000) == 32'h0);
  assign _zz_decode_IS_RS2_SIGNED = {(|_zz_decode_IS_RS2_SIGNED_5),{(|_zz_decode_IS_RS2_SIGNED_5),{(|(_zz__zz_decode_IS_RS2_SIGNED == _zz__zz_decode_IS_RS2_SIGNED_1)),{(|_zz__zz_decode_IS_RS2_SIGNED_2),{(|_zz__zz_decode_IS_RS2_SIGNED_3),{_zz__zz_decode_IS_RS2_SIGNED_4,{_zz__zz_decode_IS_RS2_SIGNED_6,_zz__zz_decode_IS_RS2_SIGNED_9}}}}}}};
  assign _zz_decode_SRC1_CTRL_2 = _zz_decode_IS_RS2_SIGNED[2 : 1];
  assign _zz_decode_SRC1_CTRL_1 = _zz_decode_SRC1_CTRL_2;
  assign _zz_decode_ALU_CTRL_2 = _zz_decode_IS_RS2_SIGNED[7 : 6];
  assign _zz_decode_ALU_CTRL_1 = _zz_decode_ALU_CTRL_2;
  assign _zz_decode_SRC2_CTRL_2 = _zz_decode_IS_RS2_SIGNED[9 : 8];
  assign _zz_decode_SRC2_CTRL_1 = _zz_decode_SRC2_CTRL_2;
  assign _zz_decode_ALU_BITWISE_CTRL_2 = _zz_decode_IS_RS2_SIGNED[19 : 18];
  assign _zz_decode_ALU_BITWISE_CTRL_1 = _zz_decode_ALU_BITWISE_CTRL_2;
  assign _zz_decode_SHIFT_CTRL_2 = _zz_decode_IS_RS2_SIGNED[22 : 21];
  assign _zz_decode_SHIFT_CTRL_1 = _zz_decode_SHIFT_CTRL_2;
  assign _zz_decode_BRANCH_CTRL_2 = _zz_decode_IS_RS2_SIGNED[24 : 23];
  assign _zz_decode_BRANCH_CTRL = _zz_decode_BRANCH_CTRL_2;
  assign _zz_decode_ENV_CTRL_2 = _zz_decode_IS_RS2_SIGNED[27 : 26];
  assign _zz_decode_ENV_CTRL_1 = _zz_decode_ENV_CTRL_2;
  assign decodeExceptionPort_valid = (decode_arbitration_isValid && (! decode_LEGAL_INSTRUCTION));
  assign decodeExceptionPort_payload_code = 4'b0010;
  assign decodeExceptionPort_payload_badAddr = decode_INSTRUCTION;
  assign when_RegFilePlugin_l63 = (decode_INSTRUCTION[11 : 7] == 5'h0);
  assign decode_RegFilePlugin_regFileReadAddress1 = decode_INSTRUCTION_ANTICIPATED[19 : 15];
  assign decode_RegFilePlugin_regFileReadAddress2 = decode_INSTRUCTION_ANTICIPATED[24 : 20];
  assign decode_RegFilePlugin_rs1Data = _zz_RegFilePlugin_regFile_port0;
  assign decode_RegFilePlugin_rs2Data = _zz_RegFilePlugin_regFile_port1;
  always @(*) begin
    lastStageRegFileWrite_valid = (_zz_lastStageRegFileWrite_valid && writeBack_arbitration_isFiring);
    if(_zz_10) begin
      lastStageRegFileWrite_valid = 1'b1;
    end
  end

  always @(*) begin
    lastStageRegFileWrite_payload_address = _zz_lastStageRegFileWrite_payload_address[11 : 7];
    if(_zz_10) begin
      lastStageRegFileWrite_payload_address = 5'h0;
    end
  end

  always @(*) begin
    lastStageRegFileWrite_payload_data = _zz_decode_RS2_2;
    if(_zz_10) begin
      lastStageRegFileWrite_payload_data = 32'h0;
    end
  end

  always @(*) begin
    case(execute_ALU_BITWISE_CTRL)
      AluBitwiseCtrlEnum_AND_1 : begin
        execute_IntAluPlugin_bitwise = (execute_SRC1 & execute_SRC2);
      end
      AluBitwiseCtrlEnum_OR_1 : begin
        execute_IntAluPlugin_bitwise = (execute_SRC1 | execute_SRC2);
      end
      default : begin
        execute_IntAluPlugin_bitwise = (execute_SRC1 ^ execute_SRC2);
      end
    endcase
  end

  always @(*) begin
    case(execute_ALU_CTRL)
      AluCtrlEnum_BITWISE : begin
        _zz_execute_REGFILE_WRITE_DATA = execute_IntAluPlugin_bitwise;
      end
      AluCtrlEnum_SLT_SLTU : begin
        _zz_execute_REGFILE_WRITE_DATA = {31'd0, _zz__zz_execute_REGFILE_WRITE_DATA};
      end
      default : begin
        _zz_execute_REGFILE_WRITE_DATA = execute_SRC_ADD_SUB;
      end
    endcase
  end

  always @(*) begin
    case(execute_SRC1_CTRL)
      Src1CtrlEnum_RS : begin
        _zz_execute_SRC1 = execute_RS1;
      end
      Src1CtrlEnum_PC_INCREMENT : begin
        _zz_execute_SRC1 = {29'd0, _zz__zz_execute_SRC1};
      end
      Src1CtrlEnum_IMU : begin
        _zz_execute_SRC1 = {execute_INSTRUCTION[31 : 12],12'h0};
      end
      default : begin
        _zz_execute_SRC1 = {27'd0, _zz__zz_execute_SRC1_1};
      end
    endcase
  end

  assign _zz_execute_SRC2_1 = execute_INSTRUCTION[31];
  always @(*) begin
    _zz_execute_SRC2_2[19] = _zz_execute_SRC2_1;
    _zz_execute_SRC2_2[18] = _zz_execute_SRC2_1;
    _zz_execute_SRC2_2[17] = _zz_execute_SRC2_1;
    _zz_execute_SRC2_2[16] = _zz_execute_SRC2_1;
    _zz_execute_SRC2_2[15] = _zz_execute_SRC2_1;
    _zz_execute_SRC2_2[14] = _zz_execute_SRC2_1;
    _zz_execute_SRC2_2[13] = _zz_execute_SRC2_1;
    _zz_execute_SRC2_2[12] = _zz_execute_SRC2_1;
    _zz_execute_SRC2_2[11] = _zz_execute_SRC2_1;
    _zz_execute_SRC2_2[10] = _zz_execute_SRC2_1;
    _zz_execute_SRC2_2[9] = _zz_execute_SRC2_1;
    _zz_execute_SRC2_2[8] = _zz_execute_SRC2_1;
    _zz_execute_SRC2_2[7] = _zz_execute_SRC2_1;
    _zz_execute_SRC2_2[6] = _zz_execute_SRC2_1;
    _zz_execute_SRC2_2[5] = _zz_execute_SRC2_1;
    _zz_execute_SRC2_2[4] = _zz_execute_SRC2_1;
    _zz_execute_SRC2_2[3] = _zz_execute_SRC2_1;
    _zz_execute_SRC2_2[2] = _zz_execute_SRC2_1;
    _zz_execute_SRC2_2[1] = _zz_execute_SRC2_1;
    _zz_execute_SRC2_2[0] = _zz_execute_SRC2_1;
  end

  assign _zz_execute_SRC2_3 = _zz__zz_execute_SRC2_3[11];
  always @(*) begin
    _zz_execute_SRC2_4[19] = _zz_execute_SRC2_3;
    _zz_execute_SRC2_4[18] = _zz_execute_SRC2_3;
    _zz_execute_SRC2_4[17] = _zz_execute_SRC2_3;
    _zz_execute_SRC2_4[16] = _zz_execute_SRC2_3;
    _zz_execute_SRC2_4[15] = _zz_execute_SRC2_3;
    _zz_execute_SRC2_4[14] = _zz_execute_SRC2_3;
    _zz_execute_SRC2_4[13] = _zz_execute_SRC2_3;
    _zz_execute_SRC2_4[12] = _zz_execute_SRC2_3;
    _zz_execute_SRC2_4[11] = _zz_execute_SRC2_3;
    _zz_execute_SRC2_4[10] = _zz_execute_SRC2_3;
    _zz_execute_SRC2_4[9] = _zz_execute_SRC2_3;
    _zz_execute_SRC2_4[8] = _zz_execute_SRC2_3;
    _zz_execute_SRC2_4[7] = _zz_execute_SRC2_3;
    _zz_execute_SRC2_4[6] = _zz_execute_SRC2_3;
    _zz_execute_SRC2_4[5] = _zz_execute_SRC2_3;
    _zz_execute_SRC2_4[4] = _zz_execute_SRC2_3;
    _zz_execute_SRC2_4[3] = _zz_execute_SRC2_3;
    _zz_execute_SRC2_4[2] = _zz_execute_SRC2_3;
    _zz_execute_SRC2_4[1] = _zz_execute_SRC2_3;
    _zz_execute_SRC2_4[0] = _zz_execute_SRC2_3;
  end

  always @(*) begin
    case(execute_SRC2_CTRL)
      Src2CtrlEnum_RS : begin
        _zz_execute_SRC2_5 = execute_RS2;
      end
      Src2CtrlEnum_IMI : begin
        _zz_execute_SRC2_5 = {_zz_execute_SRC2_2,execute_INSTRUCTION[31 : 20]};
      end
      Src2CtrlEnum_IMS : begin
        _zz_execute_SRC2_5 = {_zz_execute_SRC2_4,{execute_INSTRUCTION[31 : 25],execute_INSTRUCTION[11 : 7]}};
      end
      default : begin
        _zz_execute_SRC2_5 = _zz_execute_SRC2;
      end
    endcase
  end

  always @(*) begin
    execute_SrcPlugin_addSub = _zz_execute_SrcPlugin_addSub;
    if(execute_SRC2_FORCE_ZERO) begin
      execute_SrcPlugin_addSub = execute_SRC1;
    end
  end

  assign execute_SrcPlugin_less = ((execute_SRC1[31] == execute_SRC2[31]) ? execute_SrcPlugin_addSub[31] : (execute_SRC_LESS_UNSIGNED ? execute_SRC2[31] : execute_SRC1[31]));
  assign execute_FullBarrelShifterPlugin_amplitude = execute_SRC2[4 : 0];
  always @(*) begin
    _zz_execute_FullBarrelShifterPlugin_reversed[0] = execute_SRC1[31];
    _zz_execute_FullBarrelShifterPlugin_reversed[1] = execute_SRC1[30];
    _zz_execute_FullBarrelShifterPlugin_reversed[2] = execute_SRC1[29];
    _zz_execute_FullBarrelShifterPlugin_reversed[3] = execute_SRC1[28];
    _zz_execute_FullBarrelShifterPlugin_reversed[4] = execute_SRC1[27];
    _zz_execute_FullBarrelShifterPlugin_reversed[5] = execute_SRC1[26];
    _zz_execute_FullBarrelShifterPlugin_reversed[6] = execute_SRC1[25];
    _zz_execute_FullBarrelShifterPlugin_reversed[7] = execute_SRC1[24];
    _zz_execute_FullBarrelShifterPlugin_reversed[8] = execute_SRC1[23];
    _zz_execute_FullBarrelShifterPlugin_reversed[9] = execute_SRC1[22];
    _zz_execute_FullBarrelShifterPlugin_reversed[10] = execute_SRC1[21];
    _zz_execute_FullBarrelShifterPlugin_reversed[11] = execute_SRC1[20];
    _zz_execute_FullBarrelShifterPlugin_reversed[12] = execute_SRC1[19];
    _zz_execute_FullBarrelShifterPlugin_reversed[13] = execute_SRC1[18];
    _zz_execute_FullBarrelShifterPlugin_reversed[14] = execute_SRC1[17];
    _zz_execute_FullBarrelShifterPlugin_reversed[15] = execute_SRC1[16];
    _zz_execute_FullBarrelShifterPlugin_reversed[16] = execute_SRC1[15];
    _zz_execute_FullBarrelShifterPlugin_reversed[17] = execute_SRC1[14];
    _zz_execute_FullBarrelShifterPlugin_reversed[18] = execute_SRC1[13];
    _zz_execute_FullBarrelShifterPlugin_reversed[19] = execute_SRC1[12];
    _zz_execute_FullBarrelShifterPlugin_reversed[20] = execute_SRC1[11];
    _zz_execute_FullBarrelShifterPlugin_reversed[21] = execute_SRC1[10];
    _zz_execute_FullBarrelShifterPlugin_reversed[22] = execute_SRC1[9];
    _zz_execute_FullBarrelShifterPlugin_reversed[23] = execute_SRC1[8];
    _zz_execute_FullBarrelShifterPlugin_reversed[24] = execute_SRC1[7];
    _zz_execute_FullBarrelShifterPlugin_reversed[25] = execute_SRC1[6];
    _zz_execute_FullBarrelShifterPlugin_reversed[26] = execute_SRC1[5];
    _zz_execute_FullBarrelShifterPlugin_reversed[27] = execute_SRC1[4];
    _zz_execute_FullBarrelShifterPlugin_reversed[28] = execute_SRC1[3];
    _zz_execute_FullBarrelShifterPlugin_reversed[29] = execute_SRC1[2];
    _zz_execute_FullBarrelShifterPlugin_reversed[30] = execute_SRC1[1];
    _zz_execute_FullBarrelShifterPlugin_reversed[31] = execute_SRC1[0];
  end

  assign execute_FullBarrelShifterPlugin_reversed = ((execute_SHIFT_CTRL == ShiftCtrlEnum_SLL_1) ? _zz_execute_FullBarrelShifterPlugin_reversed : execute_SRC1);
  always @(*) begin
    _zz_decode_RS2_3[0] = memory_SHIFT_RIGHT[31];
    _zz_decode_RS2_3[1] = memory_SHIFT_RIGHT[30];
    _zz_decode_RS2_3[2] = memory_SHIFT_RIGHT[29];
    _zz_decode_RS2_3[3] = memory_SHIFT_RIGHT[28];
    _zz_decode_RS2_3[4] = memory_SHIFT_RIGHT[27];
    _zz_decode_RS2_3[5] = memory_SHIFT_RIGHT[26];
    _zz_decode_RS2_3[6] = memory_SHIFT_RIGHT[25];
    _zz_decode_RS2_3[7] = memory_SHIFT_RIGHT[24];
    _zz_decode_RS2_3[8] = memory_SHIFT_RIGHT[23];
    _zz_decode_RS2_3[9] = memory_SHIFT_RIGHT[22];
    _zz_decode_RS2_3[10] = memory_SHIFT_RIGHT[21];
    _zz_decode_RS2_3[11] = memory_SHIFT_RIGHT[20];
    _zz_decode_RS2_3[12] = memory_SHIFT_RIGHT[19];
    _zz_decode_RS2_3[13] = memory_SHIFT_RIGHT[18];
    _zz_decode_RS2_3[14] = memory_SHIFT_RIGHT[17];
    _zz_decode_RS2_3[15] = memory_SHIFT_RIGHT[16];
    _zz_decode_RS2_3[16] = memory_SHIFT_RIGHT[15];
    _zz_decode_RS2_3[17] = memory_SHIFT_RIGHT[14];
    _zz_decode_RS2_3[18] = memory_SHIFT_RIGHT[13];
    _zz_decode_RS2_3[19] = memory_SHIFT_RIGHT[12];
    _zz_decode_RS2_3[20] = memory_SHIFT_RIGHT[11];
    _zz_decode_RS2_3[21] = memory_SHIFT_RIGHT[10];
    _zz_decode_RS2_3[22] = memory_SHIFT_RIGHT[9];
    _zz_decode_RS2_3[23] = memory_SHIFT_RIGHT[8];
    _zz_decode_RS2_3[24] = memory_SHIFT_RIGHT[7];
    _zz_decode_RS2_3[25] = memory_SHIFT_RIGHT[6];
    _zz_decode_RS2_3[26] = memory_SHIFT_RIGHT[5];
    _zz_decode_RS2_3[27] = memory_SHIFT_RIGHT[4];
    _zz_decode_RS2_3[28] = memory_SHIFT_RIGHT[3];
    _zz_decode_RS2_3[29] = memory_SHIFT_RIGHT[2];
    _zz_decode_RS2_3[30] = memory_SHIFT_RIGHT[1];
    _zz_decode_RS2_3[31] = memory_SHIFT_RIGHT[0];
  end

  always @(*) begin
    HazardSimplePlugin_src0Hazard = 1'b0;
    if(when_HazardSimplePlugin_l57) begin
      if(when_HazardSimplePlugin_l58) begin
        if(when_HazardSimplePlugin_l48) begin
          HazardSimplePlugin_src0Hazard = 1'b1;
        end
      end
    end
    if(when_HazardSimplePlugin_l57_1) begin
      if(when_HazardSimplePlugin_l58_1) begin
        if(when_HazardSimplePlugin_l48_1) begin
          HazardSimplePlugin_src0Hazard = 1'b1;
        end
      end
    end
    if(when_HazardSimplePlugin_l57_2) begin
      if(when_HazardSimplePlugin_l58_2) begin
        if(when_HazardSimplePlugin_l48_2) begin
          HazardSimplePlugin_src0Hazard = 1'b1;
        end
      end
    end
    if(when_HazardSimplePlugin_l105) begin
      HazardSimplePlugin_src0Hazard = 1'b0;
    end
  end

  always @(*) begin
    HazardSimplePlugin_src1Hazard = 1'b0;
    if(when_HazardSimplePlugin_l57) begin
      if(when_HazardSimplePlugin_l58) begin
        if(when_HazardSimplePlugin_l51) begin
          HazardSimplePlugin_src1Hazard = 1'b1;
        end
      end
    end
    if(when_HazardSimplePlugin_l57_1) begin
      if(when_HazardSimplePlugin_l58_1) begin
        if(when_HazardSimplePlugin_l51_1) begin
          HazardSimplePlugin_src1Hazard = 1'b1;
        end
      end
    end
    if(when_HazardSimplePlugin_l57_2) begin
      if(when_HazardSimplePlugin_l58_2) begin
        if(when_HazardSimplePlugin_l51_2) begin
          HazardSimplePlugin_src1Hazard = 1'b1;
        end
      end
    end
    if(when_HazardSimplePlugin_l108) begin
      HazardSimplePlugin_src1Hazard = 1'b0;
    end
  end

  assign HazardSimplePlugin_writeBackWrites_valid = (_zz_lastStageRegFileWrite_valid && writeBack_arbitration_isFiring);
  assign HazardSimplePlugin_writeBackWrites_payload_address = _zz_lastStageRegFileWrite_payload_address[11 : 7];
  assign HazardSimplePlugin_writeBackWrites_payload_data = _zz_decode_RS2_2;
  assign HazardSimplePlugin_addr0Match = (HazardSimplePlugin_writeBackBuffer_payload_address == decode_INSTRUCTION[19 : 15]);
  assign HazardSimplePlugin_addr1Match = (HazardSimplePlugin_writeBackBuffer_payload_address == decode_INSTRUCTION[24 : 20]);
  assign when_HazardSimplePlugin_l47 = 1'b1;
  assign when_HazardSimplePlugin_l48 = (writeBack_INSTRUCTION[11 : 7] == decode_INSTRUCTION[19 : 15]);
  assign when_HazardSimplePlugin_l51 = (writeBack_INSTRUCTION[11 : 7] == decode_INSTRUCTION[24 : 20]);
  assign when_HazardSimplePlugin_l45 = (writeBack_arbitration_isValid && writeBack_REGFILE_WRITE_VALID);
  assign when_HazardSimplePlugin_l57 = (writeBack_arbitration_isValid && writeBack_REGFILE_WRITE_VALID);
  assign when_HazardSimplePlugin_l58 = (1'b0 || (! when_HazardSimplePlugin_l47));
  assign when_HazardSimplePlugin_l48_1 = (memory_INSTRUCTION[11 : 7] == decode_INSTRUCTION[19 : 15]);
  assign when_HazardSimplePlugin_l51_1 = (memory_INSTRUCTION[11 : 7] == decode_INSTRUCTION[24 : 20]);
  assign when_HazardSimplePlugin_l45_1 = (memory_arbitration_isValid && memory_REGFILE_WRITE_VALID);
  assign when_HazardSimplePlugin_l57_1 = (memory_arbitration_isValid && memory_REGFILE_WRITE_VALID);
  assign when_HazardSimplePlugin_l58_1 = (1'b0 || (! memory_BYPASSABLE_MEMORY_STAGE));
  assign when_HazardSimplePlugin_l48_2 = (execute_INSTRUCTION[11 : 7] == decode_INSTRUCTION[19 : 15]);
  assign when_HazardSimplePlugin_l51_2 = (execute_INSTRUCTION[11 : 7] == decode_INSTRUCTION[24 : 20]);
  assign when_HazardSimplePlugin_l45_2 = (execute_arbitration_isValid && execute_REGFILE_WRITE_VALID);
  assign when_HazardSimplePlugin_l57_2 = (execute_arbitration_isValid && execute_REGFILE_WRITE_VALID);
  assign when_HazardSimplePlugin_l58_2 = (1'b0 || (! execute_BYPASSABLE_EXECUTE_STAGE));
  assign when_HazardSimplePlugin_l105 = (! decode_RS1_USE);
  assign when_HazardSimplePlugin_l108 = (! decode_RS2_USE);
  assign when_HazardSimplePlugin_l113 = (decode_arbitration_isValid && (HazardSimplePlugin_src0Hazard || HazardSimplePlugin_src1Hazard));
  assign execute_BranchPlugin_eq = (execute_SRC1 == execute_SRC2);
  assign switch_Misc_l210_1 = execute_INSTRUCTION[14 : 12];
  always @(*) begin
    casez(switch_Misc_l210_1)
      3'b000 : begin
        _zz_execute_BRANCH_COND_RESULT = execute_BranchPlugin_eq;
      end
      3'b001 : begin
        _zz_execute_BRANCH_COND_RESULT = (! execute_BranchPlugin_eq);
      end
      3'b1?1 : begin
        _zz_execute_BRANCH_COND_RESULT = (! execute_SRC_LESS);
      end
      default : begin
        _zz_execute_BRANCH_COND_RESULT = execute_SRC_LESS;
      end
    endcase
  end

  always @(*) begin
    case(execute_BRANCH_CTRL)
      BranchCtrlEnum_INC : begin
        _zz_execute_BRANCH_COND_RESULT_1 = 1'b0;
      end
      BranchCtrlEnum_JAL : begin
        _zz_execute_BRANCH_COND_RESULT_1 = 1'b1;
      end
      BranchCtrlEnum_JALR : begin
        _zz_execute_BRANCH_COND_RESULT_1 = 1'b1;
      end
      default : begin
        _zz_execute_BRANCH_COND_RESULT_1 = _zz_execute_BRANCH_COND_RESULT;
      end
    endcase
  end

  assign _zz_execute_BranchPlugin_missAlignedTarget = execute_INSTRUCTION[31];
  always @(*) begin
    _zz_execute_BranchPlugin_missAlignedTarget_1[19] = _zz_execute_BranchPlugin_missAlignedTarget;
    _zz_execute_BranchPlugin_missAlignedTarget_1[18] = _zz_execute_BranchPlugin_missAlignedTarget;
    _zz_execute_BranchPlugin_missAlignedTarget_1[17] = _zz_execute_BranchPlugin_missAlignedTarget;
    _zz_execute_BranchPlugin_missAlignedTarget_1[16] = _zz_execute_BranchPlugin_missAlignedTarget;
    _zz_execute_BranchPlugin_missAlignedTarget_1[15] = _zz_execute_BranchPlugin_missAlignedTarget;
    _zz_execute_BranchPlugin_missAlignedTarget_1[14] = _zz_execute_BranchPlugin_missAlignedTarget;
    _zz_execute_BranchPlugin_missAlignedTarget_1[13] = _zz_execute_BranchPlugin_missAlignedTarget;
    _zz_execute_BranchPlugin_missAlignedTarget_1[12] = _zz_execute_BranchPlugin_missAlignedTarget;
    _zz_execute_BranchPlugin_missAlignedTarget_1[11] = _zz_execute_BranchPlugin_missAlignedTarget;
    _zz_execute_BranchPlugin_missAlignedTarget_1[10] = _zz_execute_BranchPlugin_missAlignedTarget;
    _zz_execute_BranchPlugin_missAlignedTarget_1[9] = _zz_execute_BranchPlugin_missAlignedTarget;
    _zz_execute_BranchPlugin_missAlignedTarget_1[8] = _zz_execute_BranchPlugin_missAlignedTarget;
    _zz_execute_BranchPlugin_missAlignedTarget_1[7] = _zz_execute_BranchPlugin_missAlignedTarget;
    _zz_execute_BranchPlugin_missAlignedTarget_1[6] = _zz_execute_BranchPlugin_missAlignedTarget;
    _zz_execute_BranchPlugin_missAlignedTarget_1[5] = _zz_execute_BranchPlugin_missAlignedTarget;
    _zz_execute_BranchPlugin_missAlignedTarget_1[4] = _zz_execute_BranchPlugin_missAlignedTarget;
    _zz_execute_BranchPlugin_missAlignedTarget_1[3] = _zz_execute_BranchPlugin_missAlignedTarget;
    _zz_execute_BranchPlugin_missAlignedTarget_1[2] = _zz_execute_BranchPlugin_missAlignedTarget;
    _zz_execute_BranchPlugin_missAlignedTarget_1[1] = _zz_execute_BranchPlugin_missAlignedTarget;
    _zz_execute_BranchPlugin_missAlignedTarget_1[0] = _zz_execute_BranchPlugin_missAlignedTarget;
  end

  assign _zz_execute_BranchPlugin_missAlignedTarget_2 = _zz__zz_execute_BranchPlugin_missAlignedTarget_2[19];
  always @(*) begin
    _zz_execute_BranchPlugin_missAlignedTarget_3[10] = _zz_execute_BranchPlugin_missAlignedTarget_2;
    _zz_execute_BranchPlugin_missAlignedTarget_3[9] = _zz_execute_BranchPlugin_missAlignedTarget_2;
    _zz_execute_BranchPlugin_missAlignedTarget_3[8] = _zz_execute_BranchPlugin_missAlignedTarget_2;
    _zz_execute_BranchPlugin_missAlignedTarget_3[7] = _zz_execute_BranchPlugin_missAlignedTarget_2;
    _zz_execute_BranchPlugin_missAlignedTarget_3[6] = _zz_execute_BranchPlugin_missAlignedTarget_2;
    _zz_execute_BranchPlugin_missAlignedTarget_3[5] = _zz_execute_BranchPlugin_missAlignedTarget_2;
    _zz_execute_BranchPlugin_missAlignedTarget_3[4] = _zz_execute_BranchPlugin_missAlignedTarget_2;
    _zz_execute_BranchPlugin_missAlignedTarget_3[3] = _zz_execute_BranchPlugin_missAlignedTarget_2;
    _zz_execute_BranchPlugin_missAlignedTarget_3[2] = _zz_execute_BranchPlugin_missAlignedTarget_2;
    _zz_execute_BranchPlugin_missAlignedTarget_3[1] = _zz_execute_BranchPlugin_missAlignedTarget_2;
    _zz_execute_BranchPlugin_missAlignedTarget_3[0] = _zz_execute_BranchPlugin_missAlignedTarget_2;
  end

  assign _zz_execute_BranchPlugin_missAlignedTarget_4 = _zz__zz_execute_BranchPlugin_missAlignedTarget_4[11];
  always @(*) begin
    _zz_execute_BranchPlugin_missAlignedTarget_5[18] = _zz_execute_BranchPlugin_missAlignedTarget_4;
    _zz_execute_BranchPlugin_missAlignedTarget_5[17] = _zz_execute_BranchPlugin_missAlignedTarget_4;
    _zz_execute_BranchPlugin_missAlignedTarget_5[16] = _zz_execute_BranchPlugin_missAlignedTarget_4;
    _zz_execute_BranchPlugin_missAlignedTarget_5[15] = _zz_execute_BranchPlugin_missAlignedTarget_4;
    _zz_execute_BranchPlugin_missAlignedTarget_5[14] = _zz_execute_BranchPlugin_missAlignedTarget_4;
    _zz_execute_BranchPlugin_missAlignedTarget_5[13] = _zz_execute_BranchPlugin_missAlignedTarget_4;
    _zz_execute_BranchPlugin_missAlignedTarget_5[12] = _zz_execute_BranchPlugin_missAlignedTarget_4;
    _zz_execute_BranchPlugin_missAlignedTarget_5[11] = _zz_execute_BranchPlugin_missAlignedTarget_4;
    _zz_execute_BranchPlugin_missAlignedTarget_5[10] = _zz_execute_BranchPlugin_missAlignedTarget_4;
    _zz_execute_BranchPlugin_missAlignedTarget_5[9] = _zz_execute_BranchPlugin_missAlignedTarget_4;
    _zz_execute_BranchPlugin_missAlignedTarget_5[8] = _zz_execute_BranchPlugin_missAlignedTarget_4;
    _zz_execute_BranchPlugin_missAlignedTarget_5[7] = _zz_execute_BranchPlugin_missAlignedTarget_4;
    _zz_execute_BranchPlugin_missAlignedTarget_5[6] = _zz_execute_BranchPlugin_missAlignedTarget_4;
    _zz_execute_BranchPlugin_missAlignedTarget_5[5] = _zz_execute_BranchPlugin_missAlignedTarget_4;
    _zz_execute_BranchPlugin_missAlignedTarget_5[4] = _zz_execute_BranchPlugin_missAlignedTarget_4;
    _zz_execute_BranchPlugin_missAlignedTarget_5[3] = _zz_execute_BranchPlugin_missAlignedTarget_4;
    _zz_execute_BranchPlugin_missAlignedTarget_5[2] = _zz_execute_BranchPlugin_missAlignedTarget_4;
    _zz_execute_BranchPlugin_missAlignedTarget_5[1] = _zz_execute_BranchPlugin_missAlignedTarget_4;
    _zz_execute_BranchPlugin_missAlignedTarget_5[0] = _zz_execute_BranchPlugin_missAlignedTarget_4;
  end

  always @(*) begin
    case(execute_BRANCH_CTRL)
      BranchCtrlEnum_JALR : begin
        _zz_execute_BranchPlugin_missAlignedTarget_6 = (_zz__zz_execute_BranchPlugin_missAlignedTarget_6[1] ^ execute_RS1[1]);
      end
      BranchCtrlEnum_JAL : begin
        _zz_execute_BranchPlugin_missAlignedTarget_6 = _zz__zz_execute_BranchPlugin_missAlignedTarget_6_1[1];
      end
      default : begin
        _zz_execute_BranchPlugin_missAlignedTarget_6 = _zz__zz_execute_BranchPlugin_missAlignedTarget_6_2[1];
      end
    endcase
  end

  assign execute_BranchPlugin_missAlignedTarget = (execute_BRANCH_COND_RESULT && _zz_execute_BranchPlugin_missAlignedTarget_6);
  always @(*) begin
    case(execute_BRANCH_CTRL)
      BranchCtrlEnum_JALR : begin
        execute_BranchPlugin_branch_src1 = execute_RS1;
      end
      default : begin
        execute_BranchPlugin_branch_src1 = execute_PC;
      end
    endcase
  end

  assign _zz_execute_BranchPlugin_branch_src2 = execute_INSTRUCTION[31];
  always @(*) begin
    _zz_execute_BranchPlugin_branch_src2_1[19] = _zz_execute_BranchPlugin_branch_src2;
    _zz_execute_BranchPlugin_branch_src2_1[18] = _zz_execute_BranchPlugin_branch_src2;
    _zz_execute_BranchPlugin_branch_src2_1[17] = _zz_execute_BranchPlugin_branch_src2;
    _zz_execute_BranchPlugin_branch_src2_1[16] = _zz_execute_BranchPlugin_branch_src2;
    _zz_execute_BranchPlugin_branch_src2_1[15] = _zz_execute_BranchPlugin_branch_src2;
    _zz_execute_BranchPlugin_branch_src2_1[14] = _zz_execute_BranchPlugin_branch_src2;
    _zz_execute_BranchPlugin_branch_src2_1[13] = _zz_execute_BranchPlugin_branch_src2;
    _zz_execute_BranchPlugin_branch_src2_1[12] = _zz_execute_BranchPlugin_branch_src2;
    _zz_execute_BranchPlugin_branch_src2_1[11] = _zz_execute_BranchPlugin_branch_src2;
    _zz_execute_BranchPlugin_branch_src2_1[10] = _zz_execute_BranchPlugin_branch_src2;
    _zz_execute_BranchPlugin_branch_src2_1[9] = _zz_execute_BranchPlugin_branch_src2;
    _zz_execute_BranchPlugin_branch_src2_1[8] = _zz_execute_BranchPlugin_branch_src2;
    _zz_execute_BranchPlugin_branch_src2_1[7] = _zz_execute_BranchPlugin_branch_src2;
    _zz_execute_BranchPlugin_branch_src2_1[6] = _zz_execute_BranchPlugin_branch_src2;
    _zz_execute_BranchPlugin_branch_src2_1[5] = _zz_execute_BranchPlugin_branch_src2;
    _zz_execute_BranchPlugin_branch_src2_1[4] = _zz_execute_BranchPlugin_branch_src2;
    _zz_execute_BranchPlugin_branch_src2_1[3] = _zz_execute_BranchPlugin_branch_src2;
    _zz_execute_BranchPlugin_branch_src2_1[2] = _zz_execute_BranchPlugin_branch_src2;
    _zz_execute_BranchPlugin_branch_src2_1[1] = _zz_execute_BranchPlugin_branch_src2;
    _zz_execute_BranchPlugin_branch_src2_1[0] = _zz_execute_BranchPlugin_branch_src2;
  end

  always @(*) begin
    case(execute_BRANCH_CTRL)
      BranchCtrlEnum_JALR : begin
        execute_BranchPlugin_branch_src2 = {_zz_execute_BranchPlugin_branch_src2_1,execute_INSTRUCTION[31 : 20]};
      end
      default : begin
        execute_BranchPlugin_branch_src2 = ((execute_BRANCH_CTRL == BranchCtrlEnum_JAL) ? {{_zz_execute_BranchPlugin_branch_src2_3,{{{_zz_execute_BranchPlugin_branch_src2_6,execute_INSTRUCTION[19 : 12]},execute_INSTRUCTION[20]},execute_INSTRUCTION[30 : 21]}},1'b0} : {{_zz_execute_BranchPlugin_branch_src2_5,{{{_zz_execute_BranchPlugin_branch_src2_7,_zz_execute_BranchPlugin_branch_src2_8},execute_INSTRUCTION[30 : 25]},execute_INSTRUCTION[11 : 8]}},1'b0});
        if(execute_PREDICTION_HAD_BRANCHED2) begin
          execute_BranchPlugin_branch_src2 = {29'd0, _zz_execute_BranchPlugin_branch_src2_9};
        end
      end
    endcase
  end

  assign _zz_execute_BranchPlugin_branch_src2_2 = _zz__zz_execute_BranchPlugin_branch_src2_2[19];
  always @(*) begin
    _zz_execute_BranchPlugin_branch_src2_3[10] = _zz_execute_BranchPlugin_branch_src2_2;
    _zz_execute_BranchPlugin_branch_src2_3[9] = _zz_execute_BranchPlugin_branch_src2_2;
    _zz_execute_BranchPlugin_branch_src2_3[8] = _zz_execute_BranchPlugin_branch_src2_2;
    _zz_execute_BranchPlugin_branch_src2_3[7] = _zz_execute_BranchPlugin_branch_src2_2;
    _zz_execute_BranchPlugin_branch_src2_3[6] = _zz_execute_BranchPlugin_branch_src2_2;
    _zz_execute_BranchPlugin_branch_src2_3[5] = _zz_execute_BranchPlugin_branch_src2_2;
    _zz_execute_BranchPlugin_branch_src2_3[4] = _zz_execute_BranchPlugin_branch_src2_2;
    _zz_execute_BranchPlugin_branch_src2_3[3] = _zz_execute_BranchPlugin_branch_src2_2;
    _zz_execute_BranchPlugin_branch_src2_3[2] = _zz_execute_BranchPlugin_branch_src2_2;
    _zz_execute_BranchPlugin_branch_src2_3[1] = _zz_execute_BranchPlugin_branch_src2_2;
    _zz_execute_BranchPlugin_branch_src2_3[0] = _zz_execute_BranchPlugin_branch_src2_2;
  end

  assign _zz_execute_BranchPlugin_branch_src2_4 = _zz__zz_execute_BranchPlugin_branch_src2_4[11];
  always @(*) begin
    _zz_execute_BranchPlugin_branch_src2_5[18] = _zz_execute_BranchPlugin_branch_src2_4;
    _zz_execute_BranchPlugin_branch_src2_5[17] = _zz_execute_BranchPlugin_branch_src2_4;
    _zz_execute_BranchPlugin_branch_src2_5[16] = _zz_execute_BranchPlugin_branch_src2_4;
    _zz_execute_BranchPlugin_branch_src2_5[15] = _zz_execute_BranchPlugin_branch_src2_4;
    _zz_execute_BranchPlugin_branch_src2_5[14] = _zz_execute_BranchPlugin_branch_src2_4;
    _zz_execute_BranchPlugin_branch_src2_5[13] = _zz_execute_BranchPlugin_branch_src2_4;
    _zz_execute_BranchPlugin_branch_src2_5[12] = _zz_execute_BranchPlugin_branch_src2_4;
    _zz_execute_BranchPlugin_branch_src2_5[11] = _zz_execute_BranchPlugin_branch_src2_4;
    _zz_execute_BranchPlugin_branch_src2_5[10] = _zz_execute_BranchPlugin_branch_src2_4;
    _zz_execute_BranchPlugin_branch_src2_5[9] = _zz_execute_BranchPlugin_branch_src2_4;
    _zz_execute_BranchPlugin_branch_src2_5[8] = _zz_execute_BranchPlugin_branch_src2_4;
    _zz_execute_BranchPlugin_branch_src2_5[7] = _zz_execute_BranchPlugin_branch_src2_4;
    _zz_execute_BranchPlugin_branch_src2_5[6] = _zz_execute_BranchPlugin_branch_src2_4;
    _zz_execute_BranchPlugin_branch_src2_5[5] = _zz_execute_BranchPlugin_branch_src2_4;
    _zz_execute_BranchPlugin_branch_src2_5[4] = _zz_execute_BranchPlugin_branch_src2_4;
    _zz_execute_BranchPlugin_branch_src2_5[3] = _zz_execute_BranchPlugin_branch_src2_4;
    _zz_execute_BranchPlugin_branch_src2_5[2] = _zz_execute_BranchPlugin_branch_src2_4;
    _zz_execute_BranchPlugin_branch_src2_5[1] = _zz_execute_BranchPlugin_branch_src2_4;
    _zz_execute_BranchPlugin_branch_src2_5[0] = _zz_execute_BranchPlugin_branch_src2_4;
  end

  assign execute_BranchPlugin_branchAdder = (execute_BranchPlugin_branch_src1 + execute_BranchPlugin_branch_src2);
  assign BranchPlugin_jumpInterface_valid = ((memory_arbitration_isValid && memory_BRANCH_DO) && (! 1'b0));
  assign BranchPlugin_jumpInterface_payload = memory_BRANCH_CALC;
  assign BranchPlugin_branchExceptionPort_valid = (memory_arbitration_isValid && (memory_BRANCH_DO && memory_BRANCH_CALC[1]));
  assign BranchPlugin_branchExceptionPort_payload_code = 4'b0000;
  assign BranchPlugin_branchExceptionPort_payload_badAddr = memory_BRANCH_CALC;
  assign IBusCachedPlugin_decodePrediction_rsp_wasWrong = BranchPlugin_jumpInterface_valid;
  always @(*) begin
    CsrPlugin_privilege = _zz_CsrPlugin_privilege;
    if(CsrPlugin_forceMachineWire) begin
      CsrPlugin_privilege = 2'b11;
    end
  end

  assign _zz_when_CsrPlugin_l965 = (CsrPlugin_mip_MTIP && CsrPlugin_mie_MTIE);
  assign _zz_when_CsrPlugin_l965_1 = (CsrPlugin_mip_MSIP && CsrPlugin_mie_MSIE);
  assign _zz_when_CsrPlugin_l965_2 = (CsrPlugin_mip_MEIP && CsrPlugin_mie_MEIE);
  assign CsrPlugin_exceptionPortCtrl_exceptionTargetPrivilegeUncapped = 2'b11;
  assign CsrPlugin_exceptionPortCtrl_exceptionTargetPrivilege = ((CsrPlugin_privilege < CsrPlugin_exceptionPortCtrl_exceptionTargetPrivilegeUncapped) ? CsrPlugin_exceptionPortCtrl_exceptionTargetPrivilegeUncapped : CsrPlugin_privilege);
  assign _zz_CsrPlugin_exceptionPortCtrl_exceptionContext_code = {decodeExceptionPort_valid,IBusCachedPlugin_decodeExceptionPort_valid};
  assign _zz_CsrPlugin_exceptionPortCtrl_exceptionContext_code_1 = _zz__zz_CsrPlugin_exceptionPortCtrl_exceptionContext_code_1[0];
  always @(*) begin
    CsrPlugin_exceptionPortCtrl_exceptionValids_decode = CsrPlugin_exceptionPortCtrl_exceptionValidsRegs_decode;
    if(_zz_when) begin
      CsrPlugin_exceptionPortCtrl_exceptionValids_decode = 1'b1;
    end
    if(decode_arbitration_isFlushed) begin
      CsrPlugin_exceptionPortCtrl_exceptionValids_decode = 1'b0;
    end
  end

  always @(*) begin
    CsrPlugin_exceptionPortCtrl_exceptionValids_execute = CsrPlugin_exceptionPortCtrl_exceptionValidsRegs_execute;
    if(CsrPlugin_selfException_valid) begin
      CsrPlugin_exceptionPortCtrl_exceptionValids_execute = 1'b1;
    end
    if(execute_arbitration_isFlushed) begin
      CsrPlugin_exceptionPortCtrl_exceptionValids_execute = 1'b0;
    end
  end

  always @(*) begin
    CsrPlugin_exceptionPortCtrl_exceptionValids_memory = CsrPlugin_exceptionPortCtrl_exceptionValidsRegs_memory;
    if(BranchPlugin_branchExceptionPort_valid) begin
      CsrPlugin_exceptionPortCtrl_exceptionValids_memory = 1'b1;
    end
    if(memory_arbitration_isFlushed) begin
      CsrPlugin_exceptionPortCtrl_exceptionValids_memory = 1'b0;
    end
  end

  always @(*) begin
    CsrPlugin_exceptionPortCtrl_exceptionValids_writeBack = CsrPlugin_exceptionPortCtrl_exceptionValidsRegs_writeBack;
    if(DBusCachedPlugin_exceptionBus_valid) begin
      CsrPlugin_exceptionPortCtrl_exceptionValids_writeBack = 1'b1;
    end
    if(writeBack_arbitration_isFlushed) begin
      CsrPlugin_exceptionPortCtrl_exceptionValids_writeBack = 1'b0;
    end
  end

  assign when_CsrPlugin_l922 = (! decode_arbitration_isStuck);
  assign when_CsrPlugin_l922_1 = (! execute_arbitration_isStuck);
  assign when_CsrPlugin_l922_2 = (! memory_arbitration_isStuck);
  assign when_CsrPlugin_l922_3 = (! writeBack_arbitration_isStuck);
  assign when_CsrPlugin_l935 = ({CsrPlugin_exceptionPortCtrl_exceptionValids_writeBack,{CsrPlugin_exceptionPortCtrl_exceptionValids_memory,{CsrPlugin_exceptionPortCtrl_exceptionValids_execute,CsrPlugin_exceptionPortCtrl_exceptionValids_decode}}} != 4'b0000);
  assign CsrPlugin_exceptionPendings_0 = CsrPlugin_exceptionPortCtrl_exceptionValidsRegs_decode;
  assign CsrPlugin_exceptionPendings_1 = CsrPlugin_exceptionPortCtrl_exceptionValidsRegs_execute;
  assign CsrPlugin_exceptionPendings_2 = CsrPlugin_exceptionPortCtrl_exceptionValidsRegs_memory;
  assign CsrPlugin_exceptionPendings_3 = CsrPlugin_exceptionPortCtrl_exceptionValidsRegs_writeBack;
  assign when_CsrPlugin_l959 = (CsrPlugin_mstatus_MIE || (CsrPlugin_privilege < 2'b11));
  assign when_CsrPlugin_l965 = ((_zz_when_CsrPlugin_l965 && 1'b1) && (! 1'b0));
  assign when_CsrPlugin_l965_1 = ((_zz_when_CsrPlugin_l965_1 && 1'b1) && (! 1'b0));
  assign when_CsrPlugin_l965_2 = ((_zz_when_CsrPlugin_l965_2 && 1'b1) && (! 1'b0));
  assign CsrPlugin_exception = (CsrPlugin_exceptionPortCtrl_exceptionValids_writeBack && CsrPlugin_allowException);
  assign CsrPlugin_pipelineLiberator_active = ((CsrPlugin_interrupt_valid && CsrPlugin_allowInterrupts) && decode_arbitration_isValid);
  assign when_CsrPlugin_l993 = (! execute_arbitration_isStuck);
  assign when_CsrPlugin_l993_1 = (! memory_arbitration_isStuck);
  assign when_CsrPlugin_l993_2 = (! writeBack_arbitration_isStuck);
  assign when_CsrPlugin_l998 = ((! CsrPlugin_pipelineLiberator_active) || decode_arbitration_removeIt);
  always @(*) begin
    CsrPlugin_pipelineLiberator_done = CsrPlugin_pipelineLiberator_pcValids_2;
    if(when_CsrPlugin_l1004) begin
      CsrPlugin_pipelineLiberator_done = 1'b0;
    end
    if(CsrPlugin_hadException) begin
      CsrPlugin_pipelineLiberator_done = 1'b0;
    end
  end

  assign when_CsrPlugin_l1004 = ({CsrPlugin_exceptionPortCtrl_exceptionValidsRegs_writeBack,{CsrPlugin_exceptionPortCtrl_exceptionValidsRegs_memory,CsrPlugin_exceptionPortCtrl_exceptionValidsRegs_execute}} != 3'b000);
  assign CsrPlugin_interruptJump = ((CsrPlugin_interrupt_valid && CsrPlugin_pipelineLiberator_done) && CsrPlugin_allowInterrupts);
  always @(*) begin
    CsrPlugin_targetPrivilege = CsrPlugin_interrupt_targetPrivilege;
    if(CsrPlugin_hadException) begin
      CsrPlugin_targetPrivilege = CsrPlugin_exceptionPortCtrl_exceptionTargetPrivilege;
    end
  end

  always @(*) begin
    CsrPlugin_trapCause = CsrPlugin_interrupt_code;
    if(CsrPlugin_hadException) begin
      CsrPlugin_trapCause = CsrPlugin_exceptionPortCtrl_exceptionContext_code;
    end
  end

  always @(*) begin
    CsrPlugin_xtvec_mode = 2'bxx;
    case(CsrPlugin_targetPrivilege)
      2'b11 : begin
        CsrPlugin_xtvec_mode = CsrPlugin_mtvec_mode;
      end
      default : begin
      end
    endcase
  end

  always @(*) begin
    CsrPlugin_xtvec_base = 30'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
    case(CsrPlugin_targetPrivilege)
      2'b11 : begin
        CsrPlugin_xtvec_base = CsrPlugin_mtvec_base;
      end
      default : begin
      end
    endcase
  end

  assign when_CsrPlugin_l1032 = (CsrPlugin_hadException || CsrPlugin_interruptJump);
  assign when_CsrPlugin_l1077 = (writeBack_arbitration_isValid && (writeBack_ENV_CTRL == EnvCtrlEnum_XRET));
  assign switch_CsrPlugin_l1081 = writeBack_INSTRUCTION[29 : 28];
  assign contextSwitching = CsrPlugin_jumpInterface_valid;
  assign when_CsrPlugin_l1121 = (execute_arbitration_isValid && (execute_ENV_CTRL == EnvCtrlEnum_WFI));
  assign when_CsrPlugin_l1123 = (! execute_CsrPlugin_wfiWake);
  assign when_CsrPlugin_l1129 = (|{(writeBack_arbitration_isValid && (writeBack_ENV_CTRL == EnvCtrlEnum_XRET)),{(memory_arbitration_isValid && (memory_ENV_CTRL == EnvCtrlEnum_XRET)),(execute_arbitration_isValid && (execute_ENV_CTRL == EnvCtrlEnum_XRET))}});
  assign execute_CsrPlugin_blockedBySideEffects = ((|{writeBack_arbitration_isValid,memory_arbitration_isValid}) || 1'b0);
  always @(*) begin
    execute_CsrPlugin_illegalAccess = 1'b1;
    if(execute_CsrPlugin_csr_3264) begin
      if(execute_CSR_READ_OPCODE) begin
        execute_CsrPlugin_illegalAccess = 1'b0;
      end
    end
    if(execute_CsrPlugin_csr_3857) begin
      if(execute_CSR_READ_OPCODE) begin
        execute_CsrPlugin_illegalAccess = 1'b0;
      end
    end
    if(execute_CsrPlugin_csr_3858) begin
      if(execute_CSR_READ_OPCODE) begin
        execute_CsrPlugin_illegalAccess = 1'b0;
      end
    end
    if(execute_CsrPlugin_csr_3859) begin
      if(execute_CSR_READ_OPCODE) begin
        execute_CsrPlugin_illegalAccess = 1'b0;
      end
    end
    if(execute_CsrPlugin_csr_3860) begin
      if(execute_CSR_READ_OPCODE) begin
        execute_CsrPlugin_illegalAccess = 1'b0;
      end
    end
    if(execute_CsrPlugin_csr_769) begin
      execute_CsrPlugin_illegalAccess = 1'b0;
    end
    if(execute_CsrPlugin_csr_768) begin
      execute_CsrPlugin_illegalAccess = 1'b0;
    end
    if(execute_CsrPlugin_csr_836) begin
      execute_CsrPlugin_illegalAccess = 1'b0;
    end
    if(execute_CsrPlugin_csr_772) begin
      execute_CsrPlugin_illegalAccess = 1'b0;
    end
    if(execute_CsrPlugin_csr_773) begin
      execute_CsrPlugin_illegalAccess = 1'b0;
    end
    if(execute_CsrPlugin_csr_833) begin
      execute_CsrPlugin_illegalAccess = 1'b0;
    end
    if(execute_CsrPlugin_csr_832) begin
      execute_CsrPlugin_illegalAccess = 1'b0;
    end
    if(execute_CsrPlugin_csr_834) begin
      execute_CsrPlugin_illegalAccess = 1'b0;
    end
    if(execute_CsrPlugin_csr_835) begin
      execute_CsrPlugin_illegalAccess = 1'b0;
    end
    if(execute_CsrPlugin_csr_2816) begin
      execute_CsrPlugin_illegalAccess = 1'b0;
    end
    if(execute_CsrPlugin_csr_2944) begin
      execute_CsrPlugin_illegalAccess = 1'b0;
    end
    if(execute_CsrPlugin_csr_2818) begin
      execute_CsrPlugin_illegalAccess = 1'b0;
    end
    if(execute_CsrPlugin_csr_2946) begin
      execute_CsrPlugin_illegalAccess = 1'b0;
    end
    if(execute_CsrPlugin_csr_3072) begin
      if(execute_CSR_READ_OPCODE) begin
        execute_CsrPlugin_illegalAccess = 1'b0;
      end
    end
    if(execute_CsrPlugin_csr_3200) begin
      if(execute_CSR_READ_OPCODE) begin
        execute_CsrPlugin_illegalAccess = 1'b0;
      end
    end
    if(execute_CsrPlugin_csr_3074) begin
      if(execute_CSR_READ_OPCODE) begin
        execute_CsrPlugin_illegalAccess = 1'b0;
      end
    end
    if(execute_CsrPlugin_csr_3202) begin
      if(execute_CSR_READ_OPCODE) begin
        execute_CsrPlugin_illegalAccess = 1'b0;
      end
    end
    if(execute_CsrPlugin_csr_3008) begin
      execute_CsrPlugin_illegalAccess = 1'b0;
    end
    if(execute_CsrPlugin_csr_4032) begin
      if(execute_CSR_READ_OPCODE) begin
        execute_CsrPlugin_illegalAccess = 1'b0;
      end
    end
    if(CsrPlugin_csrMapping_allowCsrSignal) begin
      execute_CsrPlugin_illegalAccess = 1'b0;
    end
    if(when_CsrPlugin_l1310) begin
      execute_CsrPlugin_illegalAccess = 1'b1;
    end
    if(when_CsrPlugin_l1315) begin
      execute_CsrPlugin_illegalAccess = 1'b0;
    end
  end

  always @(*) begin
    execute_CsrPlugin_illegalInstruction = 1'b0;
    if(when_CsrPlugin_l1149) begin
      if(when_CsrPlugin_l1150) begin
        execute_CsrPlugin_illegalInstruction = 1'b1;
      end
    end
  end

  always @(*) begin
    CsrPlugin_selfException_valid = 1'b0;
    if(when_CsrPlugin_l1142) begin
      CsrPlugin_selfException_valid = 1'b1;
    end
    if(when_CsrPlugin_l1157) begin
      CsrPlugin_selfException_valid = 1'b1;
    end
  end

  always @(*) begin
    CsrPlugin_selfException_payload_code = 4'bxxxx;
    if(when_CsrPlugin_l1142) begin
      CsrPlugin_selfException_payload_code = 4'b0010;
    end
    if(when_CsrPlugin_l1157) begin
      case(CsrPlugin_privilege)
        2'b00 : begin
          CsrPlugin_selfException_payload_code = 4'b1000;
        end
        default : begin
          CsrPlugin_selfException_payload_code = 4'b1011;
        end
      endcase
    end
  end

  assign CsrPlugin_selfException_payload_badAddr = execute_INSTRUCTION;
  assign when_CsrPlugin_l1142 = (execute_CsrPlugin_illegalAccess || execute_CsrPlugin_illegalInstruction);
  assign when_CsrPlugin_l1149 = (execute_arbitration_isValid && (execute_ENV_CTRL == EnvCtrlEnum_XRET));
  assign when_CsrPlugin_l1150 = (CsrPlugin_privilege < execute_INSTRUCTION[29 : 28]);
  assign when_CsrPlugin_l1157 = (execute_arbitration_isValid && (execute_ENV_CTRL == EnvCtrlEnum_ECALL));
  always @(*) begin
    execute_CsrPlugin_writeInstruction = ((execute_arbitration_isValid && execute_IS_CSR) && execute_CSR_WRITE_OPCODE);
    if(when_CsrPlugin_l1310) begin
      execute_CsrPlugin_writeInstruction = 1'b0;
    end
  end

  always @(*) begin
    execute_CsrPlugin_readInstruction = ((execute_arbitration_isValid && execute_IS_CSR) && execute_CSR_READ_OPCODE);
    if(when_CsrPlugin_l1310) begin
      execute_CsrPlugin_readInstruction = 1'b0;
    end
  end

  assign execute_CsrPlugin_writeEnable = (execute_CsrPlugin_writeInstruction && (! execute_arbitration_isStuck));
  assign execute_CsrPlugin_readEnable = (execute_CsrPlugin_readInstruction && (! execute_arbitration_isStuck));
  assign CsrPlugin_csrMapping_hazardFree = (! execute_CsrPlugin_blockedBySideEffects);
  assign execute_CsrPlugin_readToWriteData = CsrPlugin_csrMapping_readDataSignal;
  assign switch_Misc_l210_2 = execute_INSTRUCTION[13];
  always @(*) begin
    case(switch_Misc_l210_2)
      1'b0 : begin
        _zz_CsrPlugin_csrMapping_writeDataSignal = execute_SRC1;
      end
      default : begin
        _zz_CsrPlugin_csrMapping_writeDataSignal = (execute_INSTRUCTION[12] ? (execute_CsrPlugin_readToWriteData & (~ execute_SRC1)) : (execute_CsrPlugin_readToWriteData | execute_SRC1));
      end
    endcase
  end

  assign CsrPlugin_csrMapping_writeDataSignal = _zz_CsrPlugin_csrMapping_writeDataSignal;
  assign when_CsrPlugin_l1189 = (execute_arbitration_isValid && execute_IS_CSR);
  assign when_CsrPlugin_l1193 = (execute_arbitration_isValid && (execute_IS_CSR || 1'b0));
  assign execute_CsrPlugin_csrAddress = execute_INSTRUCTION[31 : 20];
  assign execute_MulPlugin_a = execute_RS1;
  assign execute_MulPlugin_b = execute_RS2;
  assign switch_MulPlugin_l87 = execute_INSTRUCTION[13 : 12];
  always @(*) begin
    case(switch_MulPlugin_l87)
      2'b01 : begin
        execute_MulPlugin_aSigned = 1'b1;
      end
      2'b10 : begin
        execute_MulPlugin_aSigned = 1'b1;
      end
      default : begin
        execute_MulPlugin_aSigned = 1'b0;
      end
    endcase
  end

  always @(*) begin
    case(switch_MulPlugin_l87)
      2'b01 : begin
        execute_MulPlugin_bSigned = 1'b1;
      end
      2'b10 : begin
        execute_MulPlugin_bSigned = 1'b0;
      end
      default : begin
        execute_MulPlugin_bSigned = 1'b0;
      end
    endcase
  end

  assign execute_MulPlugin_aULow = execute_MulPlugin_a[15 : 0];
  assign execute_MulPlugin_bULow = execute_MulPlugin_b[15 : 0];
  assign execute_MulPlugin_aSLow = {1'b0,execute_MulPlugin_a[15 : 0]};
  assign execute_MulPlugin_bSLow = {1'b0,execute_MulPlugin_b[15 : 0]};
  assign execute_MulPlugin_aHigh = {(execute_MulPlugin_aSigned && execute_MulPlugin_a[31]),execute_MulPlugin_a[31 : 16]};
  assign execute_MulPlugin_bHigh = {(execute_MulPlugin_bSigned && execute_MulPlugin_b[31]),execute_MulPlugin_b[31 : 16]};
  assign writeBack_MulPlugin_result = ($signed(_zz_writeBack_MulPlugin_result) + $signed(_zz_writeBack_MulPlugin_result_1));
  assign when_MulPlugin_l147 = (writeBack_arbitration_isValid && writeBack_IS_MUL);
  assign switch_MulPlugin_l148 = writeBack_INSTRUCTION[13 : 12];
  assign memory_DivPlugin_frontendOk = 1'b1;
  always @(*) begin
    memory_DivPlugin_div_counter_willIncrement = 1'b0;
    if(when_MulDivIterativePlugin_l128) begin
      if(when_MulDivIterativePlugin_l132) begin
        memory_DivPlugin_div_counter_willIncrement = 1'b1;
      end
    end
  end

  always @(*) begin
    memory_DivPlugin_div_counter_willClear = 1'b0;
    if(when_MulDivIterativePlugin_l162) begin
      memory_DivPlugin_div_counter_willClear = 1'b1;
    end
  end

  assign memory_DivPlugin_div_counter_willOverflowIfInc = (memory_DivPlugin_div_counter_value == 6'h21);
  assign memory_DivPlugin_div_counter_willOverflow = (memory_DivPlugin_div_counter_willOverflowIfInc && memory_DivPlugin_div_counter_willIncrement);
  always @(*) begin
    if(memory_DivPlugin_div_counter_willOverflow) begin
      memory_DivPlugin_div_counter_valueNext = 6'h0;
    end else begin
      memory_DivPlugin_div_counter_valueNext = (memory_DivPlugin_div_counter_value + _zz_memory_DivPlugin_div_counter_valueNext);
    end
    if(memory_DivPlugin_div_counter_willClear) begin
      memory_DivPlugin_div_counter_valueNext = 6'h0;
    end
  end

  assign when_MulDivIterativePlugin_l126 = (memory_DivPlugin_div_counter_value == 6'h20);
  assign when_MulDivIterativePlugin_l126_1 = (! memory_arbitration_isStuck);
  assign when_MulDivIterativePlugin_l128 = (memory_arbitration_isValid && memory_IS_DIV);
  assign when_MulDivIterativePlugin_l129 = ((! memory_DivPlugin_frontendOk) || (! memory_DivPlugin_div_done));
  assign when_MulDivIterativePlugin_l132 = (memory_DivPlugin_frontendOk && (! memory_DivPlugin_div_done));
  assign _zz_memory_DivPlugin_div_stage_0_remainderShifted = memory_DivPlugin_rs1[31 : 0];
  assign memory_DivPlugin_div_stage_0_remainderShifted = {memory_DivPlugin_accumulator[31 : 0],_zz_memory_DivPlugin_div_stage_0_remainderShifted[31]};
  assign memory_DivPlugin_div_stage_0_remainderMinusDenominator = (memory_DivPlugin_div_stage_0_remainderShifted - _zz_memory_DivPlugin_div_stage_0_remainderMinusDenominator);
  assign memory_DivPlugin_div_stage_0_outRemainder = ((! memory_DivPlugin_div_stage_0_remainderMinusDenominator[32]) ? _zz_memory_DivPlugin_div_stage_0_outRemainder : _zz_memory_DivPlugin_div_stage_0_outRemainder_1);
  assign memory_DivPlugin_div_stage_0_outNumerator = _zz_memory_DivPlugin_div_stage_0_outNumerator[31:0];
  assign when_MulDivIterativePlugin_l151 = (memory_DivPlugin_div_counter_value == 6'h20);
  assign _zz_memory_DivPlugin_div_result = (memory_INSTRUCTION[13] ? memory_DivPlugin_accumulator[31 : 0] : memory_DivPlugin_rs1[31 : 0]);
  assign when_MulDivIterativePlugin_l162 = (! memory_arbitration_isStuck);
  assign _zz_memory_DivPlugin_rs2 = (execute_RS2[31] && execute_IS_RS2_SIGNED);
  assign _zz_memory_DivPlugin_rs1 = (1'b0 || ((execute_IS_DIV && execute_RS1[31]) && execute_IS_RS1_SIGNED));
  always @(*) begin
    _zz_memory_DivPlugin_rs1_1[32] = (execute_IS_RS1_SIGNED && execute_RS1[31]);
    _zz_memory_DivPlugin_rs1_1[31 : 0] = execute_RS1;
  end

  assign _zz_CsrPlugin_csrMapping_readDataInit_1 = (_zz_CsrPlugin_csrMapping_readDataInit & externalInterruptArray_regNext);
  assign externalInterrupt = (|_zz_CsrPlugin_csrMapping_readDataInit_1);
  assign when_Pipeline_l124 = (! execute_arbitration_isStuck);
  assign when_Pipeline_l124_1 = (! memory_arbitration_isStuck);
  assign when_Pipeline_l124_2 = ((! writeBack_arbitration_isStuck) && (! CsrPlugin_exceptionPortCtrl_exceptionValids_writeBack));
  assign when_Pipeline_l124_3 = (! execute_arbitration_isStuck);
  assign when_Pipeline_l124_4 = (! memory_arbitration_isStuck);
  assign when_Pipeline_l124_5 = (! writeBack_arbitration_isStuck);
  assign when_Pipeline_l124_6 = (! execute_arbitration_isStuck);
  assign when_Pipeline_l124_7 = (! memory_arbitration_isStuck);
  assign when_Pipeline_l124_8 = (! writeBack_arbitration_isStuck);
  assign when_Pipeline_l124_9 = (! execute_arbitration_isStuck);
  assign _zz_decode_to_execute_SRC1_CTRL_1 = decode_SRC1_CTRL;
  assign _zz_decode_SRC1_CTRL = _zz_decode_SRC1_CTRL_1;
  assign when_Pipeline_l124_10 = (! execute_arbitration_isStuck);
  assign _zz_execute_SRC1_CTRL = decode_to_execute_SRC1_CTRL;
  assign when_Pipeline_l124_11 = (! execute_arbitration_isStuck);
  assign when_Pipeline_l124_12 = (! execute_arbitration_isStuck);
  assign when_Pipeline_l124_13 = (! memory_arbitration_isStuck);
  assign when_Pipeline_l124_14 = (! writeBack_arbitration_isStuck);
  assign _zz_decode_to_execute_ALU_CTRL_1 = decode_ALU_CTRL;
  assign _zz_decode_ALU_CTRL = _zz_decode_ALU_CTRL_1;
  assign when_Pipeline_l124_15 = (! execute_arbitration_isStuck);
  assign _zz_execute_ALU_CTRL = decode_to_execute_ALU_CTRL;
  assign _zz_decode_to_execute_SRC2_CTRL_1 = decode_SRC2_CTRL;
  assign _zz_decode_SRC2_CTRL = _zz_decode_SRC2_CTRL_1;
  assign when_Pipeline_l124_16 = (! execute_arbitration_isStuck);
  assign _zz_execute_SRC2_CTRL = decode_to_execute_SRC2_CTRL;
  assign when_Pipeline_l124_17 = (! execute_arbitration_isStuck);
  assign when_Pipeline_l124_18 = (! memory_arbitration_isStuck);
  assign when_Pipeline_l124_19 = (! writeBack_arbitration_isStuck);
  assign when_Pipeline_l124_20 = (! execute_arbitration_isStuck);
  assign when_Pipeline_l124_21 = (! execute_arbitration_isStuck);
  assign when_Pipeline_l124_22 = (! memory_arbitration_isStuck);
  assign when_Pipeline_l124_23 = (! execute_arbitration_isStuck);
  assign when_Pipeline_l124_24 = (! memory_arbitration_isStuck);
  assign when_Pipeline_l124_25 = (! writeBack_arbitration_isStuck);
  assign when_Pipeline_l124_26 = (! execute_arbitration_isStuck);
  assign when_Pipeline_l124_27 = (! execute_arbitration_isStuck);
  assign _zz_decode_to_execute_ALU_BITWISE_CTRL_1 = decode_ALU_BITWISE_CTRL;
  assign _zz_decode_ALU_BITWISE_CTRL = _zz_decode_ALU_BITWISE_CTRL_1;
  assign when_Pipeline_l124_28 = (! execute_arbitration_isStuck);
  assign _zz_execute_ALU_BITWISE_CTRL = decode_to_execute_ALU_BITWISE_CTRL;
  assign _zz_decode_to_execute_SHIFT_CTRL_1 = decode_SHIFT_CTRL;
  assign _zz_execute_to_memory_SHIFT_CTRL_1 = execute_SHIFT_CTRL;
  assign _zz_decode_SHIFT_CTRL = _zz_decode_SHIFT_CTRL_1;
  assign when_Pipeline_l124_29 = (! execute_arbitration_isStuck);
  assign _zz_execute_SHIFT_CTRL = decode_to_execute_SHIFT_CTRL;
  assign when_Pipeline_l124_30 = (! memory_arbitration_isStuck);
  assign _zz_memory_SHIFT_CTRL = execute_to_memory_SHIFT_CTRL;
  assign _zz_decode_to_execute_BRANCH_CTRL_1 = decode_BRANCH_CTRL;
  assign _zz_decode_BRANCH_CTRL_1 = _zz_decode_BRANCH_CTRL;
  assign when_Pipeline_l124_31 = (! execute_arbitration_isStuck);
  assign _zz_execute_BRANCH_CTRL = decode_to_execute_BRANCH_CTRL;
  assign when_Pipeline_l124_32 = (! execute_arbitration_isStuck);
  assign _zz_decode_to_execute_ENV_CTRL_1 = decode_ENV_CTRL;
  assign _zz_execute_to_memory_ENV_CTRL_1 = execute_ENV_CTRL;
  assign _zz_memory_to_writeBack_ENV_CTRL_1 = memory_ENV_CTRL;
  assign _zz_decode_ENV_CTRL = _zz_decode_ENV_CTRL_1;
  assign when_Pipeline_l124_33 = (! execute_arbitration_isStuck);
  assign _zz_execute_ENV_CTRL = decode_to_execute_ENV_CTRL;
  assign when_Pipeline_l124_34 = (! memory_arbitration_isStuck);
  assign _zz_memory_ENV_CTRL = execute_to_memory_ENV_CTRL;
  assign when_Pipeline_l124_35 = (! writeBack_arbitration_isStuck);
  assign _zz_writeBack_ENV_CTRL = memory_to_writeBack_ENV_CTRL;
  assign when_Pipeline_l124_36 = (! execute_arbitration_isStuck);
  assign when_Pipeline_l124_37 = (! memory_arbitration_isStuck);
  assign when_Pipeline_l124_38 = (! writeBack_arbitration_isStuck);
  assign when_Pipeline_l124_39 = (! execute_arbitration_isStuck);
  assign when_Pipeline_l124_40 = (! memory_arbitration_isStuck);
  assign when_Pipeline_l124_41 = (! execute_arbitration_isStuck);
  assign when_Pipeline_l124_42 = (! execute_arbitration_isStuck);
  assign when_Pipeline_l124_43 = (! execute_arbitration_isStuck);
  assign when_Pipeline_l124_44 = (! execute_arbitration_isStuck);
  assign when_Pipeline_l124_45 = (! execute_arbitration_isStuck);
  assign when_Pipeline_l124_46 = (! execute_arbitration_isStuck);
  assign when_Pipeline_l124_47 = (! execute_arbitration_isStuck);
  assign when_Pipeline_l124_48 = (! execute_arbitration_isStuck);
  assign when_Pipeline_l124_49 = (! memory_arbitration_isStuck);
  assign when_Pipeline_l124_50 = (! writeBack_arbitration_isStuck);
  assign when_Pipeline_l124_51 = (! memory_arbitration_isStuck);
  assign when_Pipeline_l124_52 = (! writeBack_arbitration_isStuck);
  assign when_Pipeline_l124_53 = (! memory_arbitration_isStuck);
  assign when_Pipeline_l124_54 = (! memory_arbitration_isStuck);
  assign when_Pipeline_l124_55 = (! memory_arbitration_isStuck);
  assign when_Pipeline_l124_56 = (! memory_arbitration_isStuck);
  assign when_Pipeline_l124_57 = (! memory_arbitration_isStuck);
  assign when_Pipeline_l124_58 = (! memory_arbitration_isStuck);
  assign when_Pipeline_l124_59 = (! memory_arbitration_isStuck);
  assign when_Pipeline_l124_60 = (! writeBack_arbitration_isStuck);
  assign when_Pipeline_l124_61 = (! writeBack_arbitration_isStuck);
  assign decode_arbitration_isFlushed = (({writeBack_arbitration_flushNext,{memory_arbitration_flushNext,execute_arbitration_flushNext}} != 3'b000) || ({writeBack_arbitration_flushIt,{memory_arbitration_flushIt,{execute_arbitration_flushIt,decode_arbitration_flushIt}}} != 4'b0000));
  assign execute_arbitration_isFlushed = (({writeBack_arbitration_flushNext,memory_arbitration_flushNext} != 2'b00) || ({writeBack_arbitration_flushIt,{memory_arbitration_flushIt,execute_arbitration_flushIt}} != 3'b000));
  assign memory_arbitration_isFlushed = ((writeBack_arbitration_flushNext != 1'b0) || ({writeBack_arbitration_flushIt,memory_arbitration_flushIt} != 2'b00));
  assign writeBack_arbitration_isFlushed = (1'b0 || (writeBack_arbitration_flushIt != 1'b0));
  assign decode_arbitration_isStuckByOthers = (decode_arbitration_haltByOther || (((1'b0 || execute_arbitration_isStuck) || memory_arbitration_isStuck) || writeBack_arbitration_isStuck));
  assign decode_arbitration_isStuck = (decode_arbitration_haltItself || decode_arbitration_isStuckByOthers);
  assign decode_arbitration_isMoving = ((! decode_arbitration_isStuck) && (! decode_arbitration_removeIt));
  assign decode_arbitration_isFiring = ((decode_arbitration_isValid && (! decode_arbitration_isStuck)) && (! decode_arbitration_removeIt));
  assign execute_arbitration_isStuckByOthers = (execute_arbitration_haltByOther || ((1'b0 || memory_arbitration_isStuck) || writeBack_arbitration_isStuck));
  assign execute_arbitration_isStuck = (execute_arbitration_haltItself || execute_arbitration_isStuckByOthers);
  assign execute_arbitration_isMoving = ((! execute_arbitration_isStuck) && (! execute_arbitration_removeIt));
  assign execute_arbitration_isFiring = ((execute_arbitration_isValid && (! execute_arbitration_isStuck)) && (! execute_arbitration_removeIt));
  assign memory_arbitration_isStuckByOthers = (memory_arbitration_haltByOther || (1'b0 || writeBack_arbitration_isStuck));
  assign memory_arbitration_isStuck = (memory_arbitration_haltItself || memory_arbitration_isStuckByOthers);
  assign memory_arbitration_isMoving = ((! memory_arbitration_isStuck) && (! memory_arbitration_removeIt));
  assign memory_arbitration_isFiring = ((memory_arbitration_isValid && (! memory_arbitration_isStuck)) && (! memory_arbitration_removeIt));
  assign writeBack_arbitration_isStuckByOthers = (writeBack_arbitration_haltByOther || 1'b0);
  assign writeBack_arbitration_isStuck = (writeBack_arbitration_haltItself || writeBack_arbitration_isStuckByOthers);
  assign writeBack_arbitration_isMoving = ((! writeBack_arbitration_isStuck) && (! writeBack_arbitration_removeIt));
  assign writeBack_arbitration_isFiring = ((writeBack_arbitration_isValid && (! writeBack_arbitration_isStuck)) && (! writeBack_arbitration_removeIt));
  assign when_Pipeline_l151 = ((! execute_arbitration_isStuck) || execute_arbitration_removeIt);
  assign when_Pipeline_l154 = ((! decode_arbitration_isStuck) && (! decode_arbitration_removeIt));
  assign when_Pipeline_l151_1 = ((! memory_arbitration_isStuck) || memory_arbitration_removeIt);
  assign when_Pipeline_l154_1 = ((! execute_arbitration_isStuck) && (! execute_arbitration_removeIt));
  assign when_Pipeline_l151_2 = ((! writeBack_arbitration_isStuck) || writeBack_arbitration_removeIt);
  assign when_Pipeline_l154_2 = ((! memory_arbitration_isStuck) && (! memory_arbitration_removeIt));
  always @(*) begin
    execute_PmpPlugin_fsm_stateNext = execute_PmpPlugin_fsm_stateReg;
    case(execute_PmpPlugin_fsm_stateReg)
      execute_PmpPlugin_fsm_enumDef_stateIdle : begin
        if(execute_PmpPlugin_fsmPending) begin
          execute_PmpPlugin_fsm_stateNext = execute_PmpPlugin_fsm_enumDef_stateWrite;
        end
      end
      execute_PmpPlugin_fsm_enumDef_stateWrite : begin
        if(execute_PmpPlugin_pmpcfgCsr_) begin
          execute_PmpPlugin_fsm_stateNext = execute_PmpPlugin_fsm_enumDef_stateCfg;
        end
        if(execute_PmpPlugin_pmpaddrCsr_) begin
          execute_PmpPlugin_fsm_stateNext = execute_PmpPlugin_fsm_enumDef_stateAddr;
        end
      end
      execute_PmpPlugin_fsm_enumDef_stateCfg : begin
        if(when_PmpPlugin_l229) begin
          execute_PmpPlugin_fsm_stateNext = execute_PmpPlugin_fsm_enumDef_stateIdle;
        end
      end
      execute_PmpPlugin_fsm_enumDef_stateAddr : begin
        execute_PmpPlugin_fsm_stateNext = execute_PmpPlugin_fsm_enumDef_stateIdle;
      end
      default : begin
      end
    endcase
    if(execute_PmpPlugin_fsm_wantStart) begin
      execute_PmpPlugin_fsm_stateNext = execute_PmpPlugin_fsm_enumDef_stateIdle;
    end
    if(execute_PmpPlugin_fsm_wantKill) begin
      execute_PmpPlugin_fsm_stateNext = execute_PmpPlugin_fsm_enumDef_BOOT;
    end
  end

  assign _zz_PmpPlugin_pmpcfg_0 = execute_PmpPlugin_writeData_[7 : 0];
  assign _zz_PmpPlugin_pmpcfg_0_1 = execute_PmpPlugin_writeData_[15 : 8];
  assign _zz_PmpPlugin_pmpcfg_0_2 = execute_PmpPlugin_writeData_[23 : 16];
  assign _zz_PmpPlugin_pmpcfg_0_3 = execute_PmpPlugin_writeData_[31 : 24];
  assign when_PmpPlugin_l209 = (! _zz_when_PmpPlugin_l209[7]);
  assign _zz_11 = ({15'd0,1'b1} <<< {execute_PmpPlugin_pmpcfgN_,2'b00});
  assign when_PmpPlugin_l209_1 = (! _zz_when_PmpPlugin_l209_1_1[7]);
  assign _zz_12 = ({15'd0,1'b1} <<< {execute_PmpPlugin_pmpcfgN_,2'b01});
  assign when_PmpPlugin_l209_2 = (! _zz_when_PmpPlugin_l209_2[7]);
  assign _zz_13 = ({15'd0,1'b1} <<< {execute_PmpPlugin_pmpcfgN_,2'b10});
  assign when_PmpPlugin_l209_3 = (! _zz_when_PmpPlugin_l209_3[7]);
  assign _zz_14 = ({15'd0,1'b1} <<< {execute_PmpPlugin_pmpcfgN_,2'b11});
  assign when_PmpPlugin_l216 = (! _zz_when_PmpPlugin_l216[7]);
  assign when_PmpPlugin_l229 = (execute_PmpPlugin_fsm_fsmCounter[1 : 0] == 2'b11);
  assign when_StateMachine_l233 = ((execute_PmpPlugin_fsm_stateReg == execute_PmpPlugin_fsm_enumDef_stateWrite) && (! (execute_PmpPlugin_fsm_stateNext == execute_PmpPlugin_fsm_enumDef_stateWrite)));
  assign when_StateMachine_l249 = ((! (execute_PmpPlugin_fsm_stateReg == execute_PmpPlugin_fsm_enumDef_stateIdle)) && (execute_PmpPlugin_fsm_stateNext == execute_PmpPlugin_fsm_enumDef_stateIdle));
  assign when_StateMachine_l249_1 = ((! (execute_PmpPlugin_fsm_stateReg == execute_PmpPlugin_fsm_enumDef_stateCfg)) && (execute_PmpPlugin_fsm_stateNext == execute_PmpPlugin_fsm_enumDef_stateCfg));
  assign when_StateMachine_l249_2 = ((! (execute_PmpPlugin_fsm_stateReg == execute_PmpPlugin_fsm_enumDef_stateAddr)) && (execute_PmpPlugin_fsm_stateNext == execute_PmpPlugin_fsm_enumDef_stateAddr));
  assign when_CsrPlugin_l1277 = (! execute_arbitration_isStuck);
  assign when_CsrPlugin_l1277_1 = (! execute_arbitration_isStuck);
  assign when_CsrPlugin_l1277_2 = (! execute_arbitration_isStuck);
  assign when_CsrPlugin_l1277_3 = (! execute_arbitration_isStuck);
  assign when_CsrPlugin_l1277_4 = (! execute_arbitration_isStuck);
  assign when_CsrPlugin_l1277_5 = (! execute_arbitration_isStuck);
  assign when_CsrPlugin_l1277_6 = (! execute_arbitration_isStuck);
  assign when_CsrPlugin_l1277_7 = (! execute_arbitration_isStuck);
  assign when_CsrPlugin_l1277_8 = (! execute_arbitration_isStuck);
  assign when_CsrPlugin_l1277_9 = (! execute_arbitration_isStuck);
  assign when_CsrPlugin_l1277_10 = (! execute_arbitration_isStuck);
  assign when_CsrPlugin_l1277_11 = (! execute_arbitration_isStuck);
  assign when_CsrPlugin_l1277_12 = (! execute_arbitration_isStuck);
  assign when_CsrPlugin_l1277_13 = (! execute_arbitration_isStuck);
  assign when_CsrPlugin_l1277_14 = (! execute_arbitration_isStuck);
  assign when_CsrPlugin_l1277_15 = (! execute_arbitration_isStuck);
  assign when_CsrPlugin_l1277_16 = (! execute_arbitration_isStuck);
  assign when_CsrPlugin_l1277_17 = (! execute_arbitration_isStuck);
  assign when_CsrPlugin_l1277_18 = (! execute_arbitration_isStuck);
  assign when_CsrPlugin_l1277_19 = (! execute_arbitration_isStuck);
  assign when_CsrPlugin_l1277_20 = (! execute_arbitration_isStuck);
  assign when_CsrPlugin_l1277_21 = (! execute_arbitration_isStuck);
  assign when_CsrPlugin_l1277_22 = (! execute_arbitration_isStuck);
  assign when_CsrPlugin_l1277_23 = (! execute_arbitration_isStuck);
  always @(*) begin
    _zz_CsrPlugin_csrMapping_readDataInit_2 = 32'h0;
    if(execute_CsrPlugin_csr_3264) begin
      _zz_CsrPlugin_csrMapping_readDataInit_2[12 : 0] = 13'h1000;
      _zz_CsrPlugin_csrMapping_readDataInit_2[25 : 20] = 6'h20;
    end
  end

  always @(*) begin
    _zz_CsrPlugin_csrMapping_readDataInit_3 = 32'h0;
    if(execute_CsrPlugin_csr_3857) begin
      _zz_CsrPlugin_csrMapping_readDataInit_3[0 : 0] = 1'b1;
    end
  end

  always @(*) begin
    _zz_CsrPlugin_csrMapping_readDataInit_4 = 32'h0;
    if(execute_CsrPlugin_csr_3858) begin
      _zz_CsrPlugin_csrMapping_readDataInit_4[1 : 0] = 2'b10;
    end
  end

  always @(*) begin
    _zz_CsrPlugin_csrMapping_readDataInit_5 = 32'h0;
    if(execute_CsrPlugin_csr_3859) begin
      _zz_CsrPlugin_csrMapping_readDataInit_5[1 : 0] = 2'b11;
    end
  end

  always @(*) begin
    _zz_CsrPlugin_csrMapping_readDataInit_6 = 32'h0;
    if(execute_CsrPlugin_csr_769) begin
      _zz_CsrPlugin_csrMapping_readDataInit_6[31 : 30] = CsrPlugin_misa_base;
      _zz_CsrPlugin_csrMapping_readDataInit_6[25 : 0] = CsrPlugin_misa_extensions;
    end
  end

  assign switch_CsrPlugin_l723 = CsrPlugin_csrMapping_writeDataSignal[12 : 11];
  always @(*) begin
    _zz_CsrPlugin_csrMapping_readDataInit_7 = 32'h0;
    if(execute_CsrPlugin_csr_768) begin
      _zz_CsrPlugin_csrMapping_readDataInit_7[7 : 7] = CsrPlugin_mstatus_MPIE;
      _zz_CsrPlugin_csrMapping_readDataInit_7[3 : 3] = CsrPlugin_mstatus_MIE;
      _zz_CsrPlugin_csrMapping_readDataInit_7[12 : 11] = CsrPlugin_mstatus_MPP;
    end
  end

  always @(*) begin
    _zz_CsrPlugin_csrMapping_readDataInit_8 = 32'h0;
    if(execute_CsrPlugin_csr_836) begin
      _zz_CsrPlugin_csrMapping_readDataInit_8[11 : 11] = CsrPlugin_mip_MEIP;
      _zz_CsrPlugin_csrMapping_readDataInit_8[7 : 7] = CsrPlugin_mip_MTIP;
      _zz_CsrPlugin_csrMapping_readDataInit_8[3 : 3] = CsrPlugin_mip_MSIP;
    end
  end

  always @(*) begin
    _zz_CsrPlugin_csrMapping_readDataInit_9 = 32'h0;
    if(execute_CsrPlugin_csr_772) begin
      _zz_CsrPlugin_csrMapping_readDataInit_9[11 : 11] = CsrPlugin_mie_MEIE;
      _zz_CsrPlugin_csrMapping_readDataInit_9[7 : 7] = CsrPlugin_mie_MTIE;
      _zz_CsrPlugin_csrMapping_readDataInit_9[3 : 3] = CsrPlugin_mie_MSIE;
    end
  end

  always @(*) begin
    _zz_CsrPlugin_csrMapping_readDataInit_10 = 32'h0;
    if(execute_CsrPlugin_csr_773) begin
      _zz_CsrPlugin_csrMapping_readDataInit_10[31 : 2] = CsrPlugin_mtvec_base;
      _zz_CsrPlugin_csrMapping_readDataInit_10[1 : 0] = CsrPlugin_mtvec_mode;
    end
  end

  always @(*) begin
    _zz_CsrPlugin_csrMapping_readDataInit_11 = 32'h0;
    if(execute_CsrPlugin_csr_833) begin
      _zz_CsrPlugin_csrMapping_readDataInit_11[31 : 0] = CsrPlugin_mepc;
    end
  end

  always @(*) begin
    _zz_CsrPlugin_csrMapping_readDataInit_12 = 32'h0;
    if(execute_CsrPlugin_csr_832) begin
      _zz_CsrPlugin_csrMapping_readDataInit_12[31 : 0] = CsrPlugin_mscratch;
    end
  end

  always @(*) begin
    _zz_CsrPlugin_csrMapping_readDataInit_13 = 32'h0;
    if(execute_CsrPlugin_csr_834) begin
      _zz_CsrPlugin_csrMapping_readDataInit_13[31 : 31] = CsrPlugin_mcause_interrupt;
      _zz_CsrPlugin_csrMapping_readDataInit_13[3 : 0] = CsrPlugin_mcause_exceptionCode;
    end
  end

  always @(*) begin
    _zz_CsrPlugin_csrMapping_readDataInit_14 = 32'h0;
    if(execute_CsrPlugin_csr_835) begin
      _zz_CsrPlugin_csrMapping_readDataInit_14[31 : 0] = CsrPlugin_mtval;
    end
  end

  always @(*) begin
    _zz_CsrPlugin_csrMapping_readDataInit_15 = 32'h0;
    if(execute_CsrPlugin_csr_2816) begin
      _zz_CsrPlugin_csrMapping_readDataInit_15[31 : 0] = CsrPlugin_mcycle[31 : 0];
    end
  end

  always @(*) begin
    _zz_CsrPlugin_csrMapping_readDataInit_16 = 32'h0;
    if(execute_CsrPlugin_csr_2944) begin
      _zz_CsrPlugin_csrMapping_readDataInit_16[31 : 0] = CsrPlugin_mcycle[63 : 32];
    end
  end

  always @(*) begin
    _zz_CsrPlugin_csrMapping_readDataInit_17 = 32'h0;
    if(execute_CsrPlugin_csr_2818) begin
      _zz_CsrPlugin_csrMapping_readDataInit_17[31 : 0] = CsrPlugin_minstret[31 : 0];
    end
  end

  always @(*) begin
    _zz_CsrPlugin_csrMapping_readDataInit_18 = 32'h0;
    if(execute_CsrPlugin_csr_2946) begin
      _zz_CsrPlugin_csrMapping_readDataInit_18[31 : 0] = CsrPlugin_minstret[63 : 32];
    end
  end

  always @(*) begin
    _zz_CsrPlugin_csrMapping_readDataInit_19 = 32'h0;
    if(execute_CsrPlugin_csr_3072) begin
      _zz_CsrPlugin_csrMapping_readDataInit_19[31 : 0] = CsrPlugin_mcycle[31 : 0];
    end
  end

  always @(*) begin
    _zz_CsrPlugin_csrMapping_readDataInit_20 = 32'h0;
    if(execute_CsrPlugin_csr_3200) begin
      _zz_CsrPlugin_csrMapping_readDataInit_20[31 : 0] = CsrPlugin_mcycle[63 : 32];
    end
  end

  always @(*) begin
    _zz_CsrPlugin_csrMapping_readDataInit_21 = 32'h0;
    if(execute_CsrPlugin_csr_3074) begin
      _zz_CsrPlugin_csrMapping_readDataInit_21[31 : 0] = CsrPlugin_minstret[31 : 0];
    end
  end

  always @(*) begin
    _zz_CsrPlugin_csrMapping_readDataInit_22 = 32'h0;
    if(execute_CsrPlugin_csr_3202) begin
      _zz_CsrPlugin_csrMapping_readDataInit_22[31 : 0] = CsrPlugin_minstret[63 : 32];
    end
  end

  always @(*) begin
    _zz_CsrPlugin_csrMapping_readDataInit_23 = 32'h0;
    if(execute_CsrPlugin_csr_3008) begin
      _zz_CsrPlugin_csrMapping_readDataInit_23[31 : 0] = _zz_CsrPlugin_csrMapping_readDataInit;
    end
  end

  always @(*) begin
    _zz_CsrPlugin_csrMapping_readDataInit_24 = 32'h0;
    if(execute_CsrPlugin_csr_4032) begin
      _zz_CsrPlugin_csrMapping_readDataInit_24[31 : 0] = _zz_CsrPlugin_csrMapping_readDataInit_1;
    end
  end

  assign CsrPlugin_csrMapping_readDataInit = (((((_zz_CsrPlugin_csrMapping_readDataInit_2 | _zz_CsrPlugin_csrMapping_readDataInit_3) | (_zz_CsrPlugin_csrMapping_readDataInit_4 | _zz_CsrPlugin_csrMapping_readDataInit_5)) | ((_zz_CsrPlugin_csrMapping_readDataInit_25 | _zz_CsrPlugin_csrMapping_readDataInit_6) | (_zz_CsrPlugin_csrMapping_readDataInit_7 | _zz_CsrPlugin_csrMapping_readDataInit_8))) | (((_zz_CsrPlugin_csrMapping_readDataInit_9 | _zz_CsrPlugin_csrMapping_readDataInit_10) | (_zz_CsrPlugin_csrMapping_readDataInit_11 | _zz_CsrPlugin_csrMapping_readDataInit_12)) | ((_zz_CsrPlugin_csrMapping_readDataInit_13 | _zz_CsrPlugin_csrMapping_readDataInit_14) | (_zz_CsrPlugin_csrMapping_readDataInit_15 | _zz_CsrPlugin_csrMapping_readDataInit_16)))) | (((_zz_CsrPlugin_csrMapping_readDataInit_17 | _zz_CsrPlugin_csrMapping_readDataInit_18) | (_zz_CsrPlugin_csrMapping_readDataInit_19 | _zz_CsrPlugin_csrMapping_readDataInit_20)) | ((_zz_CsrPlugin_csrMapping_readDataInit_21 | _zz_CsrPlugin_csrMapping_readDataInit_22) | (_zz_CsrPlugin_csrMapping_readDataInit_23 | _zz_CsrPlugin_csrMapping_readDataInit_24))));
  assign when_PmpPlugin_l155 = (CsrPlugin_privilege == 2'b11);
  assign when_PmpPlugin_l172 = ((execute_PmpPlugin_pmpcfgCsr || execute_PmpPlugin_pmpaddrCsr) && (CsrPlugin_privilege == 2'b11));
  assign when_PmpPlugin_l175 = ((! execute_PmpPlugin_fsmPending) && CsrPlugin_csrMapping_hazardFree);
  assign when_CsrPlugin_l1310 = (CsrPlugin_privilege < execute_CsrPlugin_csrAddress[9 : 8]);
  assign when_CsrPlugin_l1315 = ((! execute_arbitration_isValid) || (! execute_IS_CSR));
  assign iBusWishbone_ADR = {_zz_iBusWishbone_ADR_1,_zz_iBusWishbone_ADR};
  assign iBusWishbone_CTI = ((_zz_iBusWishbone_ADR == 3'b111) ? 3'b111 : 3'b010);
  assign iBusWishbone_BTE = 2'b00;
  assign iBusWishbone_SEL = 4'b1111;
  assign iBusWishbone_WE = 1'b0;
  assign iBusWishbone_DAT_MOSI = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
  always @(*) begin
    iBusWishbone_CYC = 1'b0;
    if(when_InstructionCache_l239) begin
      iBusWishbone_CYC = 1'b1;
    end
  end

  always @(*) begin
    iBusWishbone_STB = 1'b0;
    if(when_InstructionCache_l239) begin
      iBusWishbone_STB = 1'b1;
    end
  end

  assign when_InstructionCache_l239 = (iBus_cmd_valid || (_zz_iBusWishbone_ADR != 3'b000));
  assign iBus_cmd_ready = (iBus_cmd_valid && iBusWishbone_ACK);
  assign iBus_rsp_valid = _zz_iBus_rsp_valid;
  assign iBus_rsp_payload_data = iBusWishbone_DAT_MISO_regNext;
  assign iBus_rsp_payload_error = 1'b0;
  assign _zz_dBus_cmd_ready_5 = (dBus_cmd_payload_size == 3'b101);
  assign _zz_dBus_cmd_ready_1 = dBus_cmd_valid;
  assign _zz_dBus_cmd_ready_3 = dBus_cmd_payload_wr;
  assign _zz_dBus_cmd_ready_4 = ((! _zz_dBus_cmd_ready_5) || (_zz_dBus_cmd_ready == 3'b111));
  assign dBus_cmd_ready = (_zz_dBus_cmd_ready_2 && (_zz_dBus_cmd_ready_3 || _zz_dBus_cmd_ready_4));
  assign dBusWishbone_ADR = ((_zz_dBus_cmd_ready_5 ? {{dBus_cmd_payload_address[31 : 5],_zz_dBus_cmd_ready},2'b00} : {dBus_cmd_payload_address[31 : 2],2'b00}) >>> 2);
  assign dBusWishbone_CTI = (_zz_dBus_cmd_ready_5 ? (_zz_dBus_cmd_ready_4 ? 3'b111 : 3'b010) : 3'b000);
  assign dBusWishbone_BTE = 2'b00;
  assign dBusWishbone_SEL = (_zz_dBus_cmd_ready_3 ? dBus_cmd_payload_mask : 4'b1111);
  assign dBusWishbone_WE = _zz_dBus_cmd_ready_3;
  assign dBusWishbone_DAT_MOSI = dBus_cmd_payload_data;
  assign _zz_dBus_cmd_ready_2 = (_zz_dBus_cmd_ready_1 && dBusWishbone_ACK);
  assign dBusWishbone_CYC = _zz_dBus_cmd_ready_1;
  assign dBusWishbone_STB = _zz_dBus_cmd_ready_1;
  assign dBus_rsp_valid = _zz_dBus_rsp_valid;
  assign dBus_rsp_payload_data = dBusWishbone_DAT_MISO_regNext;
  assign dBus_rsp_payload_error = 1'b0;
  always @(posedge clk) begin
    if(reset) begin
      IBusCachedPlugin_fetchPc_pcReg <= externalResetVector;
      IBusCachedPlugin_fetchPc_correctionReg <= 1'b0;
      IBusCachedPlugin_fetchPc_booted <= 1'b0;
      IBusCachedPlugin_fetchPc_inc <= 1'b0;
      _zz_IBusCachedPlugin_iBusRsp_stages_0_output_ready_2 <= 1'b0;
      _zz_IBusCachedPlugin_iBusRsp_stages_1_output_m2sPipe_valid <= 1'b0;
      IBusCachedPlugin_injector_nextPcCalc_valids_0 <= 1'b0;
      IBusCachedPlugin_injector_nextPcCalc_valids_1 <= 1'b0;
      IBusCachedPlugin_injector_nextPcCalc_valids_2 <= 1'b0;
      IBusCachedPlugin_injector_nextPcCalc_valids_3 <= 1'b0;
      IBusCachedPlugin_injector_nextPcCalc_valids_4 <= 1'b0;
      IBusCachedPlugin_rspCounter <= 32'h0;
      dataCache_1_io_mem_cmd_rValid <= 1'b0;
      dataCache_1_io_mem_cmd_s2mPipe_rValid <= 1'b0;
      DBusCachedPlugin_rspCounter <= 32'h0;
      PmpPlugin_pmpcfg_0 <= 8'h0;
      PmpPlugin_pmpcfg_1 <= 8'h0;
      PmpPlugin_pmpcfg_2 <= 8'h0;
      PmpPlugin_pmpcfg_3 <= 8'h0;
      PmpPlugin_pmpcfg_4 <= 8'h0;
      PmpPlugin_pmpcfg_5 <= 8'h0;
      PmpPlugin_pmpcfg_6 <= 8'h0;
      PmpPlugin_pmpcfg_7 <= 8'h0;
      PmpPlugin_pmpcfg_8 <= 8'h0;
      PmpPlugin_pmpcfg_9 <= 8'h0;
      PmpPlugin_pmpcfg_10 <= 8'h0;
      PmpPlugin_pmpcfg_11 <= 8'h0;
      PmpPlugin_pmpcfg_12 <= 8'h0;
      PmpPlugin_pmpcfg_13 <= 8'h0;
      PmpPlugin_pmpcfg_14 <= 8'h0;
      PmpPlugin_pmpcfg_15 <= 8'h0;
      execute_PmpPlugin_fsmPending <= 1'b0;
      execute_PmpPlugin_pmpcfgCsr_ <= 1'b0;
      execute_PmpPlugin_pmpaddrCsr_ <= 1'b0;
      execute_PmpPlugin_fsm_fsmEnable <= 1'b0;
      execute_PmpPlugin_fsm_fsmCounter <= 4'b0000;
      _zz_10 <= 1'b1;
      HazardSimplePlugin_writeBackBuffer_valid <= 1'b0;
      _zz_CsrPlugin_privilege <= 2'b11;
      CsrPlugin_misa_base <= 2'b01;
      CsrPlugin_misa_extensions <= 26'h0101064;
      CsrPlugin_mstatus_MIE <= 1'b0;
      CsrPlugin_mstatus_MPIE <= 1'b0;
      CsrPlugin_mstatus_MPP <= 2'b11;
      CsrPlugin_mie_MEIE <= 1'b0;
      CsrPlugin_mie_MTIE <= 1'b0;
      CsrPlugin_mie_MSIE <= 1'b0;
      CsrPlugin_mcycle <= 64'h0;
      CsrPlugin_minstret <= 64'h0;
      CsrPlugin_exceptionPortCtrl_exceptionValidsRegs_decode <= 1'b0;
      CsrPlugin_exceptionPortCtrl_exceptionValidsRegs_execute <= 1'b0;
      CsrPlugin_exceptionPortCtrl_exceptionValidsRegs_memory <= 1'b0;
      CsrPlugin_exceptionPortCtrl_exceptionValidsRegs_writeBack <= 1'b0;
      CsrPlugin_interrupt_valid <= 1'b0;
      CsrPlugin_lastStageWasWfi <= 1'b0;
      CsrPlugin_pipelineLiberator_pcValids_0 <= 1'b0;
      CsrPlugin_pipelineLiberator_pcValids_1 <= 1'b0;
      CsrPlugin_pipelineLiberator_pcValids_2 <= 1'b0;
      CsrPlugin_hadException <= 1'b0;
      execute_CsrPlugin_wfiWake <= 1'b0;
      memory_DivPlugin_div_counter_value <= 6'h0;
      _zz_CsrPlugin_csrMapping_readDataInit <= 32'h0;
      execute_arbitration_isValid <= 1'b0;
      memory_arbitration_isValid <= 1'b0;
      writeBack_arbitration_isValid <= 1'b0;
      execute_PmpPlugin_fsm_stateReg <= execute_PmpPlugin_fsm_enumDef_BOOT;
      _zz_iBusWishbone_ADR <= 3'b000;
      _zz_iBus_rsp_valid <= 1'b0;
      _zz_dBus_cmd_ready <= 3'b000;
      _zz_dBus_rsp_valid <= 1'b0;
    end else begin
      if(IBusCachedPlugin_fetchPc_correction) begin
        IBusCachedPlugin_fetchPc_correctionReg <= 1'b1;
      end
      if(IBusCachedPlugin_fetchPc_output_fire) begin
        IBusCachedPlugin_fetchPc_correctionReg <= 1'b0;
      end
      IBusCachedPlugin_fetchPc_booted <= 1'b1;
      if(when_Fetcher_l134) begin
        IBusCachedPlugin_fetchPc_inc <= 1'b0;
      end
      if(IBusCachedPlugin_fetchPc_output_fire_1) begin
        IBusCachedPlugin_fetchPc_inc <= 1'b1;
      end
      if(when_Fetcher_l134_1) begin
        IBusCachedPlugin_fetchPc_inc <= 1'b0;
      end
      if(when_Fetcher_l161) begin
        IBusCachedPlugin_fetchPc_pcReg <= IBusCachedPlugin_fetchPc_pc;
      end
      if(IBusCachedPlugin_iBusRsp_flush) begin
        _zz_IBusCachedPlugin_iBusRsp_stages_0_output_ready_2 <= 1'b0;
      end
      if(_zz_IBusCachedPlugin_iBusRsp_stages_0_output_ready) begin
        _zz_IBusCachedPlugin_iBusRsp_stages_0_output_ready_2 <= (IBusCachedPlugin_iBusRsp_stages_0_output_valid && (! 1'b0));
      end
      if(IBusCachedPlugin_iBusRsp_flush) begin
        _zz_IBusCachedPlugin_iBusRsp_stages_1_output_m2sPipe_valid <= 1'b0;
      end
      if(IBusCachedPlugin_iBusRsp_stages_1_output_ready) begin
        _zz_IBusCachedPlugin_iBusRsp_stages_1_output_m2sPipe_valid <= (IBusCachedPlugin_iBusRsp_stages_1_output_valid && (! IBusCachedPlugin_iBusRsp_flush));
      end
      if(IBusCachedPlugin_fetchPc_flushed) begin
        IBusCachedPlugin_injector_nextPcCalc_valids_0 <= 1'b0;
      end
      if(when_Fetcher_l332) begin
        IBusCachedPlugin_injector_nextPcCalc_valids_0 <= 1'b1;
      end
      if(IBusCachedPlugin_fetchPc_flushed) begin
        IBusCachedPlugin_injector_nextPcCalc_valids_1 <= 1'b0;
      end
      if(when_Fetcher_l332_1) begin
        IBusCachedPlugin_injector_nextPcCalc_valids_1 <= IBusCachedPlugin_injector_nextPcCalc_valids_0;
      end
      if(IBusCachedPlugin_fetchPc_flushed) begin
        IBusCachedPlugin_injector_nextPcCalc_valids_1 <= 1'b0;
      end
      if(IBusCachedPlugin_fetchPc_flushed) begin
        IBusCachedPlugin_injector_nextPcCalc_valids_2 <= 1'b0;
      end
      if(when_Fetcher_l332_2) begin
        IBusCachedPlugin_injector_nextPcCalc_valids_2 <= IBusCachedPlugin_injector_nextPcCalc_valids_1;
      end
      if(IBusCachedPlugin_fetchPc_flushed) begin
        IBusCachedPlugin_injector_nextPcCalc_valids_2 <= 1'b0;
      end
      if(IBusCachedPlugin_fetchPc_flushed) begin
        IBusCachedPlugin_injector_nextPcCalc_valids_3 <= 1'b0;
      end
      if(when_Fetcher_l332_3) begin
        IBusCachedPlugin_injector_nextPcCalc_valids_3 <= IBusCachedPlugin_injector_nextPcCalc_valids_2;
      end
      if(IBusCachedPlugin_fetchPc_flushed) begin
        IBusCachedPlugin_injector_nextPcCalc_valids_3 <= 1'b0;
      end
      if(IBusCachedPlugin_fetchPc_flushed) begin
        IBusCachedPlugin_injector_nextPcCalc_valids_4 <= 1'b0;
      end
      if(when_Fetcher_l332_4) begin
        IBusCachedPlugin_injector_nextPcCalc_valids_4 <= IBusCachedPlugin_injector_nextPcCalc_valids_3;
      end
      if(IBusCachedPlugin_fetchPc_flushed) begin
        IBusCachedPlugin_injector_nextPcCalc_valids_4 <= 1'b0;
      end
      if(iBus_rsp_valid) begin
        IBusCachedPlugin_rspCounter <= (IBusCachedPlugin_rspCounter + 32'h00000001);
      end
      if(dataCache_1_io_mem_cmd_valid) begin
        dataCache_1_io_mem_cmd_rValid <= 1'b1;
      end
      if(dataCache_1_io_mem_cmd_s2mPipe_ready) begin
        dataCache_1_io_mem_cmd_rValid <= 1'b0;
      end
      if(dataCache_1_io_mem_cmd_s2mPipe_ready) begin
        dataCache_1_io_mem_cmd_s2mPipe_rValid <= dataCache_1_io_mem_cmd_s2mPipe_valid;
      end
      if(dBus_rsp_valid) begin
        DBusCachedPlugin_rspCounter <= (DBusCachedPlugin_rspCounter + 32'h00000001);
      end
      if(when_PmpPlugin_l138) begin
        execute_PmpPlugin_fsmPending <= 1'b0;
      end
      _zz_10 <= 1'b0;
      HazardSimplePlugin_writeBackBuffer_valid <= HazardSimplePlugin_writeBackWrites_valid;
      CsrPlugin_mcycle <= (CsrPlugin_mcycle + 64'h0000000000000001);
      if(writeBack_arbitration_isFiring) begin
        CsrPlugin_minstret <= (CsrPlugin_minstret + 64'h0000000000000001);
      end
      if(when_CsrPlugin_l922) begin
        CsrPlugin_exceptionPortCtrl_exceptionValidsRegs_decode <= 1'b0;
      end else begin
        CsrPlugin_exceptionPortCtrl_exceptionValidsRegs_decode <= CsrPlugin_exceptionPortCtrl_exceptionValids_decode;
      end
      if(when_CsrPlugin_l922_1) begin
        CsrPlugin_exceptionPortCtrl_exceptionValidsRegs_execute <= (CsrPlugin_exceptionPortCtrl_exceptionValids_decode && (! decode_arbitration_isStuck));
      end else begin
        CsrPlugin_exceptionPortCtrl_exceptionValidsRegs_execute <= CsrPlugin_exceptionPortCtrl_exceptionValids_execute;
      end
      if(when_CsrPlugin_l922_2) begin
        CsrPlugin_exceptionPortCtrl_exceptionValidsRegs_memory <= (CsrPlugin_exceptionPortCtrl_exceptionValids_execute && (! execute_arbitration_isStuck));
      end else begin
        CsrPlugin_exceptionPortCtrl_exceptionValidsRegs_memory <= CsrPlugin_exceptionPortCtrl_exceptionValids_memory;
      end
      if(when_CsrPlugin_l922_3) begin
        CsrPlugin_exceptionPortCtrl_exceptionValidsRegs_writeBack <= (CsrPlugin_exceptionPortCtrl_exceptionValids_memory && (! memory_arbitration_isStuck));
      end else begin
        CsrPlugin_exceptionPortCtrl_exceptionValidsRegs_writeBack <= 1'b0;
      end
      CsrPlugin_interrupt_valid <= 1'b0;
      if(when_CsrPlugin_l959) begin
        if(when_CsrPlugin_l965) begin
          CsrPlugin_interrupt_valid <= 1'b1;
        end
        if(when_CsrPlugin_l965_1) begin
          CsrPlugin_interrupt_valid <= 1'b1;
        end
        if(when_CsrPlugin_l965_2) begin
          CsrPlugin_interrupt_valid <= 1'b1;
        end
      end
      CsrPlugin_lastStageWasWfi <= (writeBack_arbitration_isFiring && (writeBack_ENV_CTRL == EnvCtrlEnum_WFI));
      if(CsrPlugin_pipelineLiberator_active) begin
        if(when_CsrPlugin_l993) begin
          CsrPlugin_pipelineLiberator_pcValids_0 <= 1'b1;
        end
        if(when_CsrPlugin_l993_1) begin
          CsrPlugin_pipelineLiberator_pcValids_1 <= CsrPlugin_pipelineLiberator_pcValids_0;
        end
        if(when_CsrPlugin_l993_2) begin
          CsrPlugin_pipelineLiberator_pcValids_2 <= CsrPlugin_pipelineLiberator_pcValids_1;
        end
      end
      if(when_CsrPlugin_l998) begin
        CsrPlugin_pipelineLiberator_pcValids_0 <= 1'b0;
        CsrPlugin_pipelineLiberator_pcValids_1 <= 1'b0;
        CsrPlugin_pipelineLiberator_pcValids_2 <= 1'b0;
      end
      if(CsrPlugin_interruptJump) begin
        CsrPlugin_interrupt_valid <= 1'b0;
      end
      CsrPlugin_hadException <= CsrPlugin_exception;
      if(when_CsrPlugin_l1032) begin
        _zz_CsrPlugin_privilege <= CsrPlugin_targetPrivilege;
        case(CsrPlugin_targetPrivilege)
          2'b11 : begin
            CsrPlugin_mstatus_MIE <= 1'b0;
            CsrPlugin_mstatus_MPIE <= CsrPlugin_mstatus_MIE;
            CsrPlugin_mstatus_MPP <= CsrPlugin_privilege;
          end
          default : begin
          end
        endcase
      end
      if(when_CsrPlugin_l1077) begin
        case(switch_CsrPlugin_l1081)
          2'b11 : begin
            CsrPlugin_mstatus_MPP <= 2'b00;
            CsrPlugin_mstatus_MIE <= CsrPlugin_mstatus_MPIE;
            CsrPlugin_mstatus_MPIE <= 1'b1;
            _zz_CsrPlugin_privilege <= CsrPlugin_mstatus_MPP;
          end
          default : begin
          end
        endcase
      end
      execute_CsrPlugin_wfiWake <= (({_zz_when_CsrPlugin_l965_2,{_zz_when_CsrPlugin_l965_1,_zz_when_CsrPlugin_l965}} != 3'b000) || CsrPlugin_thirdPartyWake);
      memory_DivPlugin_div_counter_value <= memory_DivPlugin_div_counter_valueNext;
      if(when_Pipeline_l151) begin
        execute_arbitration_isValid <= 1'b0;
      end
      if(when_Pipeline_l154) begin
        execute_arbitration_isValid <= decode_arbitration_isValid;
      end
      if(when_Pipeline_l151_1) begin
        memory_arbitration_isValid <= 1'b0;
      end
      if(when_Pipeline_l154_1) begin
        memory_arbitration_isValid <= execute_arbitration_isValid;
      end
      if(when_Pipeline_l151_2) begin
        writeBack_arbitration_isValid <= 1'b0;
      end
      if(when_Pipeline_l154_2) begin
        writeBack_arbitration_isValid <= memory_arbitration_isValid;
      end
      execute_PmpPlugin_fsm_stateReg <= execute_PmpPlugin_fsm_stateNext;
      case(execute_PmpPlugin_fsm_stateReg)
        execute_PmpPlugin_fsm_enumDef_stateIdle : begin
        end
        execute_PmpPlugin_fsm_enumDef_stateWrite : begin
          if(execute_PmpPlugin_pmpcfgCsr_) begin
            if(when_PmpPlugin_l209) begin
              if(_zz_11[0]) begin
                PmpPlugin_pmpcfg_0 <= _zz_PmpPlugin_pmpcfg_0;
              end
              if(_zz_11[1]) begin
                PmpPlugin_pmpcfg_1 <= _zz_PmpPlugin_pmpcfg_0;
              end
              if(_zz_11[2]) begin
                PmpPlugin_pmpcfg_2 <= _zz_PmpPlugin_pmpcfg_0;
              end
              if(_zz_11[3]) begin
                PmpPlugin_pmpcfg_3 <= _zz_PmpPlugin_pmpcfg_0;
              end
              if(_zz_11[4]) begin
                PmpPlugin_pmpcfg_4 <= _zz_PmpPlugin_pmpcfg_0;
              end
              if(_zz_11[5]) begin
                PmpPlugin_pmpcfg_5 <= _zz_PmpPlugin_pmpcfg_0;
              end
              if(_zz_11[6]) begin
                PmpPlugin_pmpcfg_6 <= _zz_PmpPlugin_pmpcfg_0;
              end
              if(_zz_11[7]) begin
                PmpPlugin_pmpcfg_7 <= _zz_PmpPlugin_pmpcfg_0;
              end
              if(_zz_11[8]) begin
                PmpPlugin_pmpcfg_8 <= _zz_PmpPlugin_pmpcfg_0;
              end
              if(_zz_11[9]) begin
                PmpPlugin_pmpcfg_9 <= _zz_PmpPlugin_pmpcfg_0;
              end
              if(_zz_11[10]) begin
                PmpPlugin_pmpcfg_10 <= _zz_PmpPlugin_pmpcfg_0;
              end
              if(_zz_11[11]) begin
                PmpPlugin_pmpcfg_11 <= _zz_PmpPlugin_pmpcfg_0;
              end
              if(_zz_11[12]) begin
                PmpPlugin_pmpcfg_12 <= _zz_PmpPlugin_pmpcfg_0;
              end
              if(_zz_11[13]) begin
                PmpPlugin_pmpcfg_13 <= _zz_PmpPlugin_pmpcfg_0;
              end
              if(_zz_11[14]) begin
                PmpPlugin_pmpcfg_14 <= _zz_PmpPlugin_pmpcfg_0;
              end
              if(_zz_11[15]) begin
                PmpPlugin_pmpcfg_15 <= _zz_PmpPlugin_pmpcfg_0;
              end
            end
            if(when_PmpPlugin_l209_1) begin
              if(_zz_12[0]) begin
                PmpPlugin_pmpcfg_0 <= _zz_PmpPlugin_pmpcfg_0_1;
              end
              if(_zz_12[1]) begin
                PmpPlugin_pmpcfg_1 <= _zz_PmpPlugin_pmpcfg_0_1;
              end
              if(_zz_12[2]) begin
                PmpPlugin_pmpcfg_2 <= _zz_PmpPlugin_pmpcfg_0_1;
              end
              if(_zz_12[3]) begin
                PmpPlugin_pmpcfg_3 <= _zz_PmpPlugin_pmpcfg_0_1;
              end
              if(_zz_12[4]) begin
                PmpPlugin_pmpcfg_4 <= _zz_PmpPlugin_pmpcfg_0_1;
              end
              if(_zz_12[5]) begin
                PmpPlugin_pmpcfg_5 <= _zz_PmpPlugin_pmpcfg_0_1;
              end
              if(_zz_12[6]) begin
                PmpPlugin_pmpcfg_6 <= _zz_PmpPlugin_pmpcfg_0_1;
              end
              if(_zz_12[7]) begin
                PmpPlugin_pmpcfg_7 <= _zz_PmpPlugin_pmpcfg_0_1;
              end
              if(_zz_12[8]) begin
                PmpPlugin_pmpcfg_8 <= _zz_PmpPlugin_pmpcfg_0_1;
              end
              if(_zz_12[9]) begin
                PmpPlugin_pmpcfg_9 <= _zz_PmpPlugin_pmpcfg_0_1;
              end
              if(_zz_12[10]) begin
                PmpPlugin_pmpcfg_10 <= _zz_PmpPlugin_pmpcfg_0_1;
              end
              if(_zz_12[11]) begin
                PmpPlugin_pmpcfg_11 <= _zz_PmpPlugin_pmpcfg_0_1;
              end
              if(_zz_12[12]) begin
                PmpPlugin_pmpcfg_12 <= _zz_PmpPlugin_pmpcfg_0_1;
              end
              if(_zz_12[13]) begin
                PmpPlugin_pmpcfg_13 <= _zz_PmpPlugin_pmpcfg_0_1;
              end
              if(_zz_12[14]) begin
                PmpPlugin_pmpcfg_14 <= _zz_PmpPlugin_pmpcfg_0_1;
              end
              if(_zz_12[15]) begin
                PmpPlugin_pmpcfg_15 <= _zz_PmpPlugin_pmpcfg_0_1;
              end
            end
            if(when_PmpPlugin_l209_2) begin
              if(_zz_13[0]) begin
                PmpPlugin_pmpcfg_0 <= _zz_PmpPlugin_pmpcfg_0_2;
              end
              if(_zz_13[1]) begin
                PmpPlugin_pmpcfg_1 <= _zz_PmpPlugin_pmpcfg_0_2;
              end
              if(_zz_13[2]) begin
                PmpPlugin_pmpcfg_2 <= _zz_PmpPlugin_pmpcfg_0_2;
              end
              if(_zz_13[3]) begin
                PmpPlugin_pmpcfg_3 <= _zz_PmpPlugin_pmpcfg_0_2;
              end
              if(_zz_13[4]) begin
                PmpPlugin_pmpcfg_4 <= _zz_PmpPlugin_pmpcfg_0_2;
              end
              if(_zz_13[5]) begin
                PmpPlugin_pmpcfg_5 <= _zz_PmpPlugin_pmpcfg_0_2;
              end
              if(_zz_13[6]) begin
                PmpPlugin_pmpcfg_6 <= _zz_PmpPlugin_pmpcfg_0_2;
              end
              if(_zz_13[7]) begin
                PmpPlugin_pmpcfg_7 <= _zz_PmpPlugin_pmpcfg_0_2;
              end
              if(_zz_13[8]) begin
                PmpPlugin_pmpcfg_8 <= _zz_PmpPlugin_pmpcfg_0_2;
              end
              if(_zz_13[9]) begin
                PmpPlugin_pmpcfg_9 <= _zz_PmpPlugin_pmpcfg_0_2;
              end
              if(_zz_13[10]) begin
                PmpPlugin_pmpcfg_10 <= _zz_PmpPlugin_pmpcfg_0_2;
              end
              if(_zz_13[11]) begin
                PmpPlugin_pmpcfg_11 <= _zz_PmpPlugin_pmpcfg_0_2;
              end
              if(_zz_13[12]) begin
                PmpPlugin_pmpcfg_12 <= _zz_PmpPlugin_pmpcfg_0_2;
              end
              if(_zz_13[13]) begin
                PmpPlugin_pmpcfg_13 <= _zz_PmpPlugin_pmpcfg_0_2;
              end
              if(_zz_13[14]) begin
                PmpPlugin_pmpcfg_14 <= _zz_PmpPlugin_pmpcfg_0_2;
              end
              if(_zz_13[15]) begin
                PmpPlugin_pmpcfg_15 <= _zz_PmpPlugin_pmpcfg_0_2;
              end
            end
            if(when_PmpPlugin_l209_3) begin
              if(_zz_14[0]) begin
                PmpPlugin_pmpcfg_0 <= _zz_PmpPlugin_pmpcfg_0_3;
              end
              if(_zz_14[1]) begin
                PmpPlugin_pmpcfg_1 <= _zz_PmpPlugin_pmpcfg_0_3;
              end
              if(_zz_14[2]) begin
                PmpPlugin_pmpcfg_2 <= _zz_PmpPlugin_pmpcfg_0_3;
              end
              if(_zz_14[3]) begin
                PmpPlugin_pmpcfg_3 <= _zz_PmpPlugin_pmpcfg_0_3;
              end
              if(_zz_14[4]) begin
                PmpPlugin_pmpcfg_4 <= _zz_PmpPlugin_pmpcfg_0_3;
              end
              if(_zz_14[5]) begin
                PmpPlugin_pmpcfg_5 <= _zz_PmpPlugin_pmpcfg_0_3;
              end
              if(_zz_14[6]) begin
                PmpPlugin_pmpcfg_6 <= _zz_PmpPlugin_pmpcfg_0_3;
              end
              if(_zz_14[7]) begin
                PmpPlugin_pmpcfg_7 <= _zz_PmpPlugin_pmpcfg_0_3;
              end
              if(_zz_14[8]) begin
                PmpPlugin_pmpcfg_8 <= _zz_PmpPlugin_pmpcfg_0_3;
              end
              if(_zz_14[9]) begin
                PmpPlugin_pmpcfg_9 <= _zz_PmpPlugin_pmpcfg_0_3;
              end
              if(_zz_14[10]) begin
                PmpPlugin_pmpcfg_10 <= _zz_PmpPlugin_pmpcfg_0_3;
              end
              if(_zz_14[11]) begin
                PmpPlugin_pmpcfg_11 <= _zz_PmpPlugin_pmpcfg_0_3;
              end
              if(_zz_14[12]) begin
                PmpPlugin_pmpcfg_12 <= _zz_PmpPlugin_pmpcfg_0_3;
              end
              if(_zz_14[13]) begin
                PmpPlugin_pmpcfg_13 <= _zz_PmpPlugin_pmpcfg_0_3;
              end
              if(_zz_14[14]) begin
                PmpPlugin_pmpcfg_14 <= _zz_PmpPlugin_pmpcfg_0_3;
              end
              if(_zz_14[15]) begin
                PmpPlugin_pmpcfg_15 <= _zz_PmpPlugin_pmpcfg_0_3;
              end
            end
          end
        end
        execute_PmpPlugin_fsm_enumDef_stateCfg : begin
          execute_PmpPlugin_fsm_fsmCounter <= (execute_PmpPlugin_fsm_fsmCounter + 4'b0001);
        end
        execute_PmpPlugin_fsm_enumDef_stateAddr : begin
        end
        default : begin
        end
      endcase
      if(when_StateMachine_l233) begin
        execute_PmpPlugin_fsm_fsmEnable <= 1'b1;
      end
      if(when_StateMachine_l249) begin
        execute_PmpPlugin_fsmPending <= 1'b0;
        execute_PmpPlugin_fsm_fsmEnable <= 1'b0;
        execute_PmpPlugin_fsm_fsmCounter <= 4'b0000;
      end
      if(when_StateMachine_l249_1) begin
        execute_PmpPlugin_fsm_fsmCounter <= {execute_PmpPlugin_pmpcfgN_,2'b00};
      end
      if(when_StateMachine_l249_2) begin
        execute_PmpPlugin_fsm_fsmCounter <= execute_PmpPlugin_pmpNcfg_;
      end
      if(execute_CsrPlugin_csr_769) begin
        if(execute_CsrPlugin_writeEnable) begin
          CsrPlugin_misa_base <= CsrPlugin_csrMapping_writeDataSignal[31 : 30];
          CsrPlugin_misa_extensions <= CsrPlugin_csrMapping_writeDataSignal[25 : 0];
        end
      end
      if(execute_CsrPlugin_csr_768) begin
        if(execute_CsrPlugin_writeEnable) begin
          CsrPlugin_mstatus_MPIE <= CsrPlugin_csrMapping_writeDataSignal[7];
          CsrPlugin_mstatus_MIE <= CsrPlugin_csrMapping_writeDataSignal[3];
          case(switch_CsrPlugin_l723)
            2'b11 : begin
              CsrPlugin_mstatus_MPP <= 2'b11;
            end
            2'b00 : begin
              CsrPlugin_mstatus_MPP <= 2'b00;
            end
            default : begin
            end
          endcase
        end
      end
      if(execute_CsrPlugin_csr_772) begin
        if(execute_CsrPlugin_writeEnable) begin
          CsrPlugin_mie_MEIE <= CsrPlugin_csrMapping_writeDataSignal[11];
          CsrPlugin_mie_MTIE <= CsrPlugin_csrMapping_writeDataSignal[7];
          CsrPlugin_mie_MSIE <= CsrPlugin_csrMapping_writeDataSignal[3];
        end
      end
      if(execute_CsrPlugin_csr_2816) begin
        if(execute_CsrPlugin_writeEnable) begin
          CsrPlugin_mcycle[31 : 0] <= CsrPlugin_csrMapping_writeDataSignal[31 : 0];
        end
      end
      if(execute_CsrPlugin_csr_2944) begin
        if(execute_CsrPlugin_writeEnable) begin
          CsrPlugin_mcycle[63 : 32] <= CsrPlugin_csrMapping_writeDataSignal[31 : 0];
        end
      end
      if(execute_CsrPlugin_csr_2818) begin
        if(execute_CsrPlugin_writeEnable) begin
          CsrPlugin_minstret[31 : 0] <= CsrPlugin_csrMapping_writeDataSignal[31 : 0];
        end
      end
      if(execute_CsrPlugin_csr_2946) begin
        if(execute_CsrPlugin_writeEnable) begin
          CsrPlugin_minstret[63 : 32] <= CsrPlugin_csrMapping_writeDataSignal[31 : 0];
        end
      end
      if(execute_CsrPlugin_csr_3008) begin
        if(execute_CsrPlugin_writeEnable) begin
          _zz_CsrPlugin_csrMapping_readDataInit <= CsrPlugin_csrMapping_writeDataSignal[31 : 0];
        end
      end
      if(execute_CsrPlugin_writeInstruction) begin
        if(when_PmpPlugin_l172) begin
          if(when_PmpPlugin_l175) begin
            execute_PmpPlugin_fsmPending <= 1'b1;
            execute_PmpPlugin_pmpcfgCsr_ <= execute_PmpPlugin_pmpcfgCsr;
            execute_PmpPlugin_pmpaddrCsr_ <= execute_PmpPlugin_pmpaddrCsr;
          end
        end
      end
      if(when_InstructionCache_l239) begin
        if(iBusWishbone_ACK) begin
          _zz_iBusWishbone_ADR <= (_zz_iBusWishbone_ADR + 3'b001);
        end
      end
      _zz_iBus_rsp_valid <= (iBusWishbone_CYC && iBusWishbone_ACK);
      if((_zz_dBus_cmd_ready_1 && _zz_dBus_cmd_ready_2)) begin
        _zz_dBus_cmd_ready <= (_zz_dBus_cmd_ready + 3'b001);
        if(_zz_dBus_cmd_ready_4) begin
          _zz_dBus_cmd_ready <= 3'b000;
        end
      end
      _zz_dBus_rsp_valid <= ((_zz_dBus_cmd_ready_1 && (! dBusWishbone_WE)) && dBusWishbone_ACK);
    end
  end

  always @(posedge clk) begin
    if(IBusCachedPlugin_iBusRsp_stages_1_output_ready) begin
      _zz_IBusCachedPlugin_iBusRsp_stages_1_output_m2sPipe_payload <= IBusCachedPlugin_iBusRsp_stages_1_output_payload;
    end
    if(IBusCachedPlugin_iBusRsp_stages_1_input_ready) begin
      IBusCachedPlugin_s1_tightlyCoupledHit <= IBusCachedPlugin_s0_tightlyCoupledHit;
    end
    if(IBusCachedPlugin_iBusRsp_stages_2_input_ready) begin
      IBusCachedPlugin_s2_tightlyCoupledHit <= IBusCachedPlugin_s1_tightlyCoupledHit;
    end
    if(dataCache_1_io_mem_cmd_ready) begin
      dataCache_1_io_mem_cmd_rData_wr <= dataCache_1_io_mem_cmd_payload_wr;
      dataCache_1_io_mem_cmd_rData_uncached <= dataCache_1_io_mem_cmd_payload_uncached;
      dataCache_1_io_mem_cmd_rData_address <= dataCache_1_io_mem_cmd_payload_address;
      dataCache_1_io_mem_cmd_rData_data <= dataCache_1_io_mem_cmd_payload_data;
      dataCache_1_io_mem_cmd_rData_mask <= dataCache_1_io_mem_cmd_payload_mask;
      dataCache_1_io_mem_cmd_rData_size <= dataCache_1_io_mem_cmd_payload_size;
      dataCache_1_io_mem_cmd_rData_last <= dataCache_1_io_mem_cmd_payload_last;
    end
    if(dataCache_1_io_mem_cmd_s2mPipe_ready) begin
      dataCache_1_io_mem_cmd_s2mPipe_rData_wr <= dataCache_1_io_mem_cmd_s2mPipe_payload_wr;
      dataCache_1_io_mem_cmd_s2mPipe_rData_uncached <= dataCache_1_io_mem_cmd_s2mPipe_payload_uncached;
      dataCache_1_io_mem_cmd_s2mPipe_rData_address <= dataCache_1_io_mem_cmd_s2mPipe_payload_address;
      dataCache_1_io_mem_cmd_s2mPipe_rData_data <= dataCache_1_io_mem_cmd_s2mPipe_payload_data;
      dataCache_1_io_mem_cmd_s2mPipe_rData_mask <= dataCache_1_io_mem_cmd_s2mPipe_payload_mask;
      dataCache_1_io_mem_cmd_s2mPipe_rData_size <= dataCache_1_io_mem_cmd_s2mPipe_payload_size;
      dataCache_1_io_mem_cmd_s2mPipe_rData_last <= dataCache_1_io_mem_cmd_s2mPipe_payload_last;
    end
    if(when_PmpPlugin_l246) begin
      if(_zz_8[0]) begin
        PmpPlugin_base_0 <= PmpPlugin_setter_io_base;
      end
      if(_zz_8[1]) begin
        PmpPlugin_base_1 <= PmpPlugin_setter_io_base;
      end
      if(_zz_8[2]) begin
        PmpPlugin_base_2 <= PmpPlugin_setter_io_base;
      end
      if(_zz_8[3]) begin
        PmpPlugin_base_3 <= PmpPlugin_setter_io_base;
      end
      if(_zz_8[4]) begin
        PmpPlugin_base_4 <= PmpPlugin_setter_io_base;
      end
      if(_zz_8[5]) begin
        PmpPlugin_base_5 <= PmpPlugin_setter_io_base;
      end
      if(_zz_8[6]) begin
        PmpPlugin_base_6 <= PmpPlugin_setter_io_base;
      end
      if(_zz_8[7]) begin
        PmpPlugin_base_7 <= PmpPlugin_setter_io_base;
      end
      if(_zz_8[8]) begin
        PmpPlugin_base_8 <= PmpPlugin_setter_io_base;
      end
      if(_zz_8[9]) begin
        PmpPlugin_base_9 <= PmpPlugin_setter_io_base;
      end
      if(_zz_8[10]) begin
        PmpPlugin_base_10 <= PmpPlugin_setter_io_base;
      end
      if(_zz_8[11]) begin
        PmpPlugin_base_11 <= PmpPlugin_setter_io_base;
      end
      if(_zz_8[12]) begin
        PmpPlugin_base_12 <= PmpPlugin_setter_io_base;
      end
      if(_zz_8[13]) begin
        PmpPlugin_base_13 <= PmpPlugin_setter_io_base;
      end
      if(_zz_8[14]) begin
        PmpPlugin_base_14 <= PmpPlugin_setter_io_base;
      end
      if(_zz_8[15]) begin
        PmpPlugin_base_15 <= PmpPlugin_setter_io_base;
      end
      if(_zz_9[0]) begin
        PmpPlugin_mask_0 <= PmpPlugin_setter_io_mask;
      end
      if(_zz_9[1]) begin
        PmpPlugin_mask_1 <= PmpPlugin_setter_io_mask;
      end
      if(_zz_9[2]) begin
        PmpPlugin_mask_2 <= PmpPlugin_setter_io_mask;
      end
      if(_zz_9[3]) begin
        PmpPlugin_mask_3 <= PmpPlugin_setter_io_mask;
      end
      if(_zz_9[4]) begin
        PmpPlugin_mask_4 <= PmpPlugin_setter_io_mask;
      end
      if(_zz_9[5]) begin
        PmpPlugin_mask_5 <= PmpPlugin_setter_io_mask;
      end
      if(_zz_9[6]) begin
        PmpPlugin_mask_6 <= PmpPlugin_setter_io_mask;
      end
      if(_zz_9[7]) begin
        PmpPlugin_mask_7 <= PmpPlugin_setter_io_mask;
      end
      if(_zz_9[8]) begin
        PmpPlugin_mask_8 <= PmpPlugin_setter_io_mask;
      end
      if(_zz_9[9]) begin
        PmpPlugin_mask_9 <= PmpPlugin_setter_io_mask;
      end
      if(_zz_9[10]) begin
        PmpPlugin_mask_10 <= PmpPlugin_setter_io_mask;
      end
      if(_zz_9[11]) begin
        PmpPlugin_mask_11 <= PmpPlugin_setter_io_mask;
      end
      if(_zz_9[12]) begin
        PmpPlugin_mask_12 <= PmpPlugin_setter_io_mask;
      end
      if(_zz_9[13]) begin
        PmpPlugin_mask_13 <= PmpPlugin_setter_io_mask;
      end
      if(_zz_9[14]) begin
        PmpPlugin_mask_14 <= PmpPlugin_setter_io_mask;
      end
      if(_zz_9[15]) begin
        PmpPlugin_mask_15 <= PmpPlugin_setter_io_mask;
      end
    end
    HazardSimplePlugin_writeBackBuffer_payload_address <= HazardSimplePlugin_writeBackWrites_payload_address;
    HazardSimplePlugin_writeBackBuffer_payload_data <= HazardSimplePlugin_writeBackWrites_payload_data;
    CsrPlugin_mip_MEIP <= externalInterrupt;
    CsrPlugin_mip_MTIP <= timerInterrupt;
    CsrPlugin_mip_MSIP <= softwareInterrupt;
    if(_zz_when) begin
      CsrPlugin_exceptionPortCtrl_exceptionContext_code <= (_zz_CsrPlugin_exceptionPortCtrl_exceptionContext_code_1 ? IBusCachedPlugin_decodeExceptionPort_payload_code : decodeExceptionPort_payload_code);
      CsrPlugin_exceptionPortCtrl_exceptionContext_badAddr <= (_zz_CsrPlugin_exceptionPortCtrl_exceptionContext_code_1 ? IBusCachedPlugin_decodeExceptionPort_payload_badAddr : decodeExceptionPort_payload_badAddr);
    end
    if(CsrPlugin_selfException_valid) begin
      CsrPlugin_exceptionPortCtrl_exceptionContext_code <= CsrPlugin_selfException_payload_code;
      CsrPlugin_exceptionPortCtrl_exceptionContext_badAddr <= CsrPlugin_selfException_payload_badAddr;
    end
    if(BranchPlugin_branchExceptionPort_valid) begin
      CsrPlugin_exceptionPortCtrl_exceptionContext_code <= BranchPlugin_branchExceptionPort_payload_code;
      CsrPlugin_exceptionPortCtrl_exceptionContext_badAddr <= BranchPlugin_branchExceptionPort_payload_badAddr;
    end
    if(DBusCachedPlugin_exceptionBus_valid) begin
      CsrPlugin_exceptionPortCtrl_exceptionContext_code <= DBusCachedPlugin_exceptionBus_payload_code;
      CsrPlugin_exceptionPortCtrl_exceptionContext_badAddr <= DBusCachedPlugin_exceptionBus_payload_badAddr;
    end
    if(when_CsrPlugin_l959) begin
      if(when_CsrPlugin_l965) begin
        CsrPlugin_interrupt_code <= 4'b0111;
        CsrPlugin_interrupt_targetPrivilege <= 2'b11;
      end
      if(when_CsrPlugin_l965_1) begin
        CsrPlugin_interrupt_code <= 4'b0011;
        CsrPlugin_interrupt_targetPrivilege <= 2'b11;
      end
      if(when_CsrPlugin_l965_2) begin
        CsrPlugin_interrupt_code <= 4'b1011;
        CsrPlugin_interrupt_targetPrivilege <= 2'b11;
      end
    end
    if(when_CsrPlugin_l1032) begin
      case(CsrPlugin_targetPrivilege)
        2'b11 : begin
          CsrPlugin_mcause_interrupt <= (! CsrPlugin_hadException);
          CsrPlugin_mcause_exceptionCode <= CsrPlugin_trapCause;
          CsrPlugin_mepc <= writeBack_PC;
          if(CsrPlugin_hadException) begin
            CsrPlugin_mtval <= CsrPlugin_exceptionPortCtrl_exceptionContext_badAddr;
          end
        end
        default : begin
        end
      endcase
    end
    if(when_MulDivIterativePlugin_l126) begin
      memory_DivPlugin_div_done <= 1'b1;
    end
    if(when_MulDivIterativePlugin_l126_1) begin
      memory_DivPlugin_div_done <= 1'b0;
    end
    if(when_MulDivIterativePlugin_l128) begin
      if(when_MulDivIterativePlugin_l132) begin
        memory_DivPlugin_rs1[31 : 0] <= memory_DivPlugin_div_stage_0_outNumerator;
        memory_DivPlugin_accumulator[31 : 0] <= memory_DivPlugin_div_stage_0_outRemainder;
        if(when_MulDivIterativePlugin_l151) begin
          memory_DivPlugin_div_result <= _zz_memory_DivPlugin_div_result_1[31:0];
        end
      end
    end
    if(when_MulDivIterativePlugin_l162) begin
      memory_DivPlugin_accumulator <= 65'h0;
      memory_DivPlugin_rs1 <= ((_zz_memory_DivPlugin_rs1 ? (~ _zz_memory_DivPlugin_rs1_1) : _zz_memory_DivPlugin_rs1_1) + _zz_memory_DivPlugin_rs1_2);
      memory_DivPlugin_rs2 <= ((_zz_memory_DivPlugin_rs2 ? (~ execute_RS2) : execute_RS2) + _zz_memory_DivPlugin_rs2_1);
      memory_DivPlugin_div_needRevert <= ((_zz_memory_DivPlugin_rs1 ^ (_zz_memory_DivPlugin_rs2 && (! execute_INSTRUCTION[13]))) && (! (((execute_RS2 == 32'h0) && execute_IS_RS2_SIGNED) && (! execute_INSTRUCTION[13]))));
    end
    externalInterruptArray_regNext <= externalInterruptArray;
    if(when_Pipeline_l124) begin
      decode_to_execute_PC <= decode_PC;
    end
    if(when_Pipeline_l124_1) begin
      execute_to_memory_PC <= _zz_execute_SRC2;
    end
    if(when_Pipeline_l124_2) begin
      memory_to_writeBack_PC <= memory_PC;
    end
    if(when_Pipeline_l124_3) begin
      decode_to_execute_INSTRUCTION <= decode_INSTRUCTION;
    end
    if(when_Pipeline_l124_4) begin
      execute_to_memory_INSTRUCTION <= execute_INSTRUCTION;
    end
    if(when_Pipeline_l124_5) begin
      memory_to_writeBack_INSTRUCTION <= memory_INSTRUCTION;
    end
    if(when_Pipeline_l124_6) begin
      decode_to_execute_FORMAL_PC_NEXT <= _zz_decode_to_execute_FORMAL_PC_NEXT;
    end
    if(when_Pipeline_l124_7) begin
      execute_to_memory_FORMAL_PC_NEXT <= execute_FORMAL_PC_NEXT;
    end
    if(when_Pipeline_l124_8) begin
      memory_to_writeBack_FORMAL_PC_NEXT <= _zz_memory_to_writeBack_FORMAL_PC_NEXT;
    end
    if(when_Pipeline_l124_9) begin
      decode_to_execute_MEMORY_FORCE_CONSTISTENCY <= decode_MEMORY_FORCE_CONSTISTENCY;
    end
    if(when_Pipeline_l124_10) begin
      decode_to_execute_SRC1_CTRL <= _zz_decode_to_execute_SRC1_CTRL;
    end
    if(when_Pipeline_l124_11) begin
      decode_to_execute_SRC_USE_SUB_LESS <= decode_SRC_USE_SUB_LESS;
    end
    if(when_Pipeline_l124_12) begin
      decode_to_execute_MEMORY_ENABLE <= decode_MEMORY_ENABLE;
    end
    if(when_Pipeline_l124_13) begin
      execute_to_memory_MEMORY_ENABLE <= execute_MEMORY_ENABLE;
    end
    if(when_Pipeline_l124_14) begin
      memory_to_writeBack_MEMORY_ENABLE <= memory_MEMORY_ENABLE;
    end
    if(when_Pipeline_l124_15) begin
      decode_to_execute_ALU_CTRL <= _zz_decode_to_execute_ALU_CTRL;
    end
    if(when_Pipeline_l124_16) begin
      decode_to_execute_SRC2_CTRL <= _zz_decode_to_execute_SRC2_CTRL;
    end
    if(when_Pipeline_l124_17) begin
      decode_to_execute_REGFILE_WRITE_VALID <= decode_REGFILE_WRITE_VALID;
    end
    if(when_Pipeline_l124_18) begin
      execute_to_memory_REGFILE_WRITE_VALID <= execute_REGFILE_WRITE_VALID;
    end
    if(when_Pipeline_l124_19) begin
      memory_to_writeBack_REGFILE_WRITE_VALID <= memory_REGFILE_WRITE_VALID;
    end
    if(when_Pipeline_l124_20) begin
      decode_to_execute_BYPASSABLE_EXECUTE_STAGE <= decode_BYPASSABLE_EXECUTE_STAGE;
    end
    if(when_Pipeline_l124_21) begin
      decode_to_execute_BYPASSABLE_MEMORY_STAGE <= decode_BYPASSABLE_MEMORY_STAGE;
    end
    if(when_Pipeline_l124_22) begin
      execute_to_memory_BYPASSABLE_MEMORY_STAGE <= execute_BYPASSABLE_MEMORY_STAGE;
    end
    if(when_Pipeline_l124_23) begin
      decode_to_execute_MEMORY_WR <= decode_MEMORY_WR;
    end
    if(when_Pipeline_l124_24) begin
      execute_to_memory_MEMORY_WR <= execute_MEMORY_WR;
    end
    if(when_Pipeline_l124_25) begin
      memory_to_writeBack_MEMORY_WR <= memory_MEMORY_WR;
    end
    if(when_Pipeline_l124_26) begin
      decode_to_execute_MEMORY_MANAGMENT <= decode_MEMORY_MANAGMENT;
    end
    if(when_Pipeline_l124_27) begin
      decode_to_execute_SRC_LESS_UNSIGNED <= decode_SRC_LESS_UNSIGNED;
    end
    if(when_Pipeline_l124_28) begin
      decode_to_execute_ALU_BITWISE_CTRL <= _zz_decode_to_execute_ALU_BITWISE_CTRL;
    end
    if(when_Pipeline_l124_29) begin
      decode_to_execute_SHIFT_CTRL <= _zz_decode_to_execute_SHIFT_CTRL;
    end
    if(when_Pipeline_l124_30) begin
      execute_to_memory_SHIFT_CTRL <= _zz_execute_to_memory_SHIFT_CTRL;
    end
    if(when_Pipeline_l124_31) begin
      decode_to_execute_BRANCH_CTRL <= _zz_decode_to_execute_BRANCH_CTRL;
    end
    if(when_Pipeline_l124_32) begin
      decode_to_execute_IS_CSR <= decode_IS_CSR;
    end
    if(when_Pipeline_l124_33) begin
      decode_to_execute_ENV_CTRL <= _zz_decode_to_execute_ENV_CTRL;
    end
    if(when_Pipeline_l124_34) begin
      execute_to_memory_ENV_CTRL <= _zz_execute_to_memory_ENV_CTRL;
    end
    if(when_Pipeline_l124_35) begin
      memory_to_writeBack_ENV_CTRL <= _zz_memory_to_writeBack_ENV_CTRL;
    end
    if(when_Pipeline_l124_36) begin
      decode_to_execute_IS_MUL <= decode_IS_MUL;
    end
    if(when_Pipeline_l124_37) begin
      execute_to_memory_IS_MUL <= execute_IS_MUL;
    end
    if(when_Pipeline_l124_38) begin
      memory_to_writeBack_IS_MUL <= memory_IS_MUL;
    end
    if(when_Pipeline_l124_39) begin
      decode_to_execute_IS_DIV <= decode_IS_DIV;
    end
    if(when_Pipeline_l124_40) begin
      execute_to_memory_IS_DIV <= execute_IS_DIV;
    end
    if(when_Pipeline_l124_41) begin
      decode_to_execute_IS_RS1_SIGNED <= decode_IS_RS1_SIGNED;
    end
    if(when_Pipeline_l124_42) begin
      decode_to_execute_IS_RS2_SIGNED <= decode_IS_RS2_SIGNED;
    end
    if(when_Pipeline_l124_43) begin
      decode_to_execute_RS1 <= decode_RS1;
    end
    if(when_Pipeline_l124_44) begin
      decode_to_execute_RS2 <= decode_RS2;
    end
    if(when_Pipeline_l124_45) begin
      decode_to_execute_SRC2_FORCE_ZERO <= decode_SRC2_FORCE_ZERO;
    end
    if(when_Pipeline_l124_46) begin
      decode_to_execute_PREDICTION_HAD_BRANCHED2 <= decode_PREDICTION_HAD_BRANCHED2;
    end
    if(when_Pipeline_l124_47) begin
      decode_to_execute_CSR_WRITE_OPCODE <= decode_CSR_WRITE_OPCODE;
    end
    if(when_Pipeline_l124_48) begin
      decode_to_execute_CSR_READ_OPCODE <= decode_CSR_READ_OPCODE;
    end
    if(when_Pipeline_l124_49) begin
      execute_to_memory_MEMORY_STORE_DATA_RF <= execute_MEMORY_STORE_DATA_RF;
    end
    if(when_Pipeline_l124_50) begin
      memory_to_writeBack_MEMORY_STORE_DATA_RF <= memory_MEMORY_STORE_DATA_RF;
    end
    if(when_Pipeline_l124_51) begin
      execute_to_memory_REGFILE_WRITE_DATA <= _zz_decode_RS2;
    end
    if(when_Pipeline_l124_52) begin
      memory_to_writeBack_REGFILE_WRITE_DATA <= _zz_decode_RS2_1;
    end
    if(when_Pipeline_l124_53) begin
      execute_to_memory_SHIFT_RIGHT <= execute_SHIFT_RIGHT;
    end
    if(when_Pipeline_l124_54) begin
      execute_to_memory_BRANCH_DO <= execute_BRANCH_DO;
    end
    if(when_Pipeline_l124_55) begin
      execute_to_memory_BRANCH_CALC <= execute_BRANCH_CALC;
    end
    if(when_Pipeline_l124_56) begin
      execute_to_memory_MUL_LL <= execute_MUL_LL;
    end
    if(when_Pipeline_l124_57) begin
      execute_to_memory_MUL_LH <= execute_MUL_LH;
    end
    if(when_Pipeline_l124_58) begin
      execute_to_memory_MUL_HL <= execute_MUL_HL;
    end
    if(when_Pipeline_l124_59) begin
      execute_to_memory_MUL_HH <= execute_MUL_HH;
    end
    if(when_Pipeline_l124_60) begin
      memory_to_writeBack_MUL_HH <= memory_MUL_HH;
    end
    if(when_Pipeline_l124_61) begin
      memory_to_writeBack_MUL_LOW <= memory_MUL_LOW;
    end
    if(when_CsrPlugin_l1277) begin
      execute_CsrPlugin_csr_3264 <= (decode_INSTRUCTION[31 : 20] == 12'hcc0);
    end
    if(when_CsrPlugin_l1277_1) begin
      execute_CsrPlugin_csr_3857 <= (decode_INSTRUCTION[31 : 20] == 12'hf11);
    end
    if(when_CsrPlugin_l1277_2) begin
      execute_CsrPlugin_csr_3858 <= (decode_INSTRUCTION[31 : 20] == 12'hf12);
    end
    if(when_CsrPlugin_l1277_3) begin
      execute_CsrPlugin_csr_3859 <= (decode_INSTRUCTION[31 : 20] == 12'hf13);
    end
    if(when_CsrPlugin_l1277_4) begin
      execute_CsrPlugin_csr_3860 <= (decode_INSTRUCTION[31 : 20] == 12'hf14);
    end
    if(when_CsrPlugin_l1277_5) begin
      execute_CsrPlugin_csr_769 <= (decode_INSTRUCTION[31 : 20] == 12'h301);
    end
    if(when_CsrPlugin_l1277_6) begin
      execute_CsrPlugin_csr_768 <= (decode_INSTRUCTION[31 : 20] == 12'h300);
    end
    if(when_CsrPlugin_l1277_7) begin
      execute_CsrPlugin_csr_836 <= (decode_INSTRUCTION[31 : 20] == 12'h344);
    end
    if(when_CsrPlugin_l1277_8) begin
      execute_CsrPlugin_csr_772 <= (decode_INSTRUCTION[31 : 20] == 12'h304);
    end
    if(when_CsrPlugin_l1277_9) begin
      execute_CsrPlugin_csr_773 <= (decode_INSTRUCTION[31 : 20] == 12'h305);
    end
    if(when_CsrPlugin_l1277_10) begin
      execute_CsrPlugin_csr_833 <= (decode_INSTRUCTION[31 : 20] == 12'h341);
    end
    if(when_CsrPlugin_l1277_11) begin
      execute_CsrPlugin_csr_832 <= (decode_INSTRUCTION[31 : 20] == 12'h340);
    end
    if(when_CsrPlugin_l1277_12) begin
      execute_CsrPlugin_csr_834 <= (decode_INSTRUCTION[31 : 20] == 12'h342);
    end
    if(when_CsrPlugin_l1277_13) begin
      execute_CsrPlugin_csr_835 <= (decode_INSTRUCTION[31 : 20] == 12'h343);
    end
    if(when_CsrPlugin_l1277_14) begin
      execute_CsrPlugin_csr_2816 <= (decode_INSTRUCTION[31 : 20] == 12'hb00);
    end
    if(when_CsrPlugin_l1277_15) begin
      execute_CsrPlugin_csr_2944 <= (decode_INSTRUCTION[31 : 20] == 12'hb80);
    end
    if(when_CsrPlugin_l1277_16) begin
      execute_CsrPlugin_csr_2818 <= (decode_INSTRUCTION[31 : 20] == 12'hb02);
    end
    if(when_CsrPlugin_l1277_17) begin
      execute_CsrPlugin_csr_2946 <= (decode_INSTRUCTION[31 : 20] == 12'hb82);
    end
    if(when_CsrPlugin_l1277_18) begin
      execute_CsrPlugin_csr_3072 <= (decode_INSTRUCTION[31 : 20] == 12'hc00);
    end
    if(when_CsrPlugin_l1277_19) begin
      execute_CsrPlugin_csr_3200 <= (decode_INSTRUCTION[31 : 20] == 12'hc80);
    end
    if(when_CsrPlugin_l1277_20) begin
      execute_CsrPlugin_csr_3074 <= (decode_INSTRUCTION[31 : 20] == 12'hc02);
    end
    if(when_CsrPlugin_l1277_21) begin
      execute_CsrPlugin_csr_3202 <= (decode_INSTRUCTION[31 : 20] == 12'hc82);
    end
    if(when_CsrPlugin_l1277_22) begin
      execute_CsrPlugin_csr_3008 <= (decode_INSTRUCTION[31 : 20] == 12'hbc0);
    end
    if(when_CsrPlugin_l1277_23) begin
      execute_CsrPlugin_csr_4032 <= (decode_INSTRUCTION[31 : 20] == 12'hfc0);
    end
    if(execute_CsrPlugin_csr_836) begin
      if(execute_CsrPlugin_writeEnable) begin
        CsrPlugin_mip_MSIP <= CsrPlugin_csrMapping_writeDataSignal[3];
      end
    end
    if(execute_CsrPlugin_csr_773) begin
      if(execute_CsrPlugin_writeEnable) begin
        CsrPlugin_mtvec_base <= CsrPlugin_csrMapping_writeDataSignal[31 : 2];
        CsrPlugin_mtvec_mode <= CsrPlugin_csrMapping_writeDataSignal[1 : 0];
      end
    end
    if(execute_CsrPlugin_csr_833) begin
      if(execute_CsrPlugin_writeEnable) begin
        CsrPlugin_mepc <= CsrPlugin_csrMapping_writeDataSignal[31 : 0];
      end
    end
    if(execute_CsrPlugin_csr_832) begin
      if(execute_CsrPlugin_writeEnable) begin
        CsrPlugin_mscratch <= CsrPlugin_csrMapping_writeDataSignal[31 : 0];
      end
    end
    if(execute_CsrPlugin_csr_834) begin
      if(execute_CsrPlugin_writeEnable) begin
        CsrPlugin_mcause_interrupt <= CsrPlugin_csrMapping_writeDataSignal[31];
        CsrPlugin_mcause_exceptionCode <= CsrPlugin_csrMapping_writeDataSignal[3 : 0];
      end
    end
    if(execute_CsrPlugin_csr_835) begin
      if(execute_CsrPlugin_writeEnable) begin
        CsrPlugin_mtval <= CsrPlugin_csrMapping_writeDataSignal[31 : 0];
      end
    end
    if(execute_CsrPlugin_writeInstruction) begin
      if(when_PmpPlugin_l172) begin
        if(when_PmpPlugin_l175) begin
          execute_PmpPlugin_writeData_ <= CsrPlugin_csrMapping_writeDataSignal;
          execute_PmpPlugin_pmpNcfg_ <= execute_PmpPlugin_pmpNcfg;
          execute_PmpPlugin_pmpcfgN_ <= execute_PmpPlugin_pmpcfgN;
        end
      end
    end
    iBusWishbone_DAT_MISO_regNext <= iBusWishbone_DAT_MISO;
    dBusWishbone_DAT_MISO_regNext <= dBusWishbone_DAT_MISO;
  end


endmodule

module DataCache (
  input               io_cpu_execute_isValid,
  input      [31:0]   io_cpu_execute_address,
  output reg          io_cpu_execute_haltIt,
  input               io_cpu_execute_args_wr,
  input      [1:0]    io_cpu_execute_args_size,
  input               io_cpu_execute_args_totalyConsistent,
  output              io_cpu_execute_refilling,
  input               io_cpu_memory_isValid,
  input               io_cpu_memory_isStuck,
  output              io_cpu_memory_isWrite,
  input      [31:0]   io_cpu_memory_address,
  input      [31:0]   io_cpu_memory_mmuRsp_physicalAddress,
  input               io_cpu_memory_mmuRsp_isIoAccess,
  input               io_cpu_memory_mmuRsp_isPaging,
  input               io_cpu_memory_mmuRsp_allowRead,
  input               io_cpu_memory_mmuRsp_allowWrite,
  input               io_cpu_memory_mmuRsp_allowExecute,
  input               io_cpu_memory_mmuRsp_exception,
  input               io_cpu_memory_mmuRsp_refilling,
  input               io_cpu_memory_mmuRsp_bypassTranslation,
  input               io_cpu_writeBack_isValid,
  input               io_cpu_writeBack_isStuck,
  input               io_cpu_writeBack_isFiring,
  input               io_cpu_writeBack_isUser,
  output reg          io_cpu_writeBack_haltIt,
  output              io_cpu_writeBack_isWrite,
  input      [31:0]   io_cpu_writeBack_storeData,
  output reg [31:0]   io_cpu_writeBack_data,
  input      [31:0]   io_cpu_writeBack_address,
  output              io_cpu_writeBack_mmuException,
  output              io_cpu_writeBack_unalignedAccess,
  output reg          io_cpu_writeBack_accessError,
  output              io_cpu_writeBack_keepMemRspData,
  input               io_cpu_writeBack_fence_SW,
  input               io_cpu_writeBack_fence_SR,
  input               io_cpu_writeBack_fence_SO,
  input               io_cpu_writeBack_fence_SI,
  input               io_cpu_writeBack_fence_PW,
  input               io_cpu_writeBack_fence_PR,
  input               io_cpu_writeBack_fence_PO,
  input               io_cpu_writeBack_fence_PI,
  input      [3:0]    io_cpu_writeBack_fence_FM,
  output              io_cpu_writeBack_exclusiveOk,
  output reg          io_cpu_redo,
  input               io_cpu_flush_valid,
  output              io_cpu_flush_ready,
  input               io_cpu_flush_payload_singleLine,
  input      [6:0]    io_cpu_flush_payload_lineId,
  output reg          io_mem_cmd_valid,
  input               io_mem_cmd_ready,
  output reg          io_mem_cmd_payload_wr,
  output              io_mem_cmd_payload_uncached,
  output reg [31:0]   io_mem_cmd_payload_address,
  output     [31:0]   io_mem_cmd_payload_data,
  output     [3:0]    io_mem_cmd_payload_mask,
  output reg [2:0]    io_mem_cmd_payload_size,
  output              io_mem_cmd_payload_last,
  input               io_mem_rsp_valid,
  input               io_mem_rsp_payload_last,
  input      [31:0]   io_mem_rsp_payload_data,
  input               io_mem_rsp_payload_error,
  input               clk,
  input               reset
);

  reg        [21:0]   _zz_ways_0_tags_port0;
  reg        [31:0]   _zz_ways_0_data_port0;
  wire       [21:0]   _zz_ways_0_tags_port;
  wire       [9:0]    _zz_stage0_dataColisions;
  wire       [9:0]    _zz__zz_stageA_dataColisions;
  wire       [0:0]    _zz_when;
  wire       [2:0]    _zz_loader_counter_valueNext;
  wire       [0:0]    _zz_loader_counter_valueNext_1;
  wire       [1:0]    _zz_loader_waysAllocator;
  reg                 _zz_1;
  reg                 _zz_2;
  wire                haltCpu;
  reg                 tagsReadCmd_valid;
  reg        [6:0]    tagsReadCmd_payload;
  reg                 tagsWriteCmd_valid;
  reg        [0:0]    tagsWriteCmd_payload_way;
  reg        [6:0]    tagsWriteCmd_payload_address;
  reg                 tagsWriteCmd_payload_data_valid;
  reg                 tagsWriteCmd_payload_data_error;
  reg        [19:0]   tagsWriteCmd_payload_data_address;
  reg                 tagsWriteLastCmd_valid;
  reg        [0:0]    tagsWriteLastCmd_payload_way;
  reg        [6:0]    tagsWriteLastCmd_payload_address;
  reg                 tagsWriteLastCmd_payload_data_valid;
  reg                 tagsWriteLastCmd_payload_data_error;
  reg        [19:0]   tagsWriteLastCmd_payload_data_address;
  reg                 dataReadCmd_valid;
  reg        [9:0]    dataReadCmd_payload;
  reg                 dataWriteCmd_valid;
  reg        [0:0]    dataWriteCmd_payload_way;
  reg        [9:0]    dataWriteCmd_payload_address;
  reg        [31:0]   dataWriteCmd_payload_data;
  reg        [3:0]    dataWriteCmd_payload_mask;
  wire                _zz_ways_0_tagsReadRsp_valid;
  wire                ways_0_tagsReadRsp_valid;
  wire                ways_0_tagsReadRsp_error;
  wire       [19:0]   ways_0_tagsReadRsp_address;
  wire       [21:0]   _zz_ways_0_tagsReadRsp_valid_1;
  wire                _zz_ways_0_dataReadRspMem;
  wire       [31:0]   ways_0_dataReadRspMem;
  wire       [31:0]   ways_0_dataReadRsp;
  wire                when_DataCache_l642;
  wire                when_DataCache_l645;
  wire                when_DataCache_l664;
  wire                rspSync;
  wire                rspLast;
  reg                 memCmdSent;
  wire                io_mem_cmd_fire;
  wire                when_DataCache_l686;
  reg        [3:0]    _zz_stage0_mask;
  wire       [3:0]    stage0_mask;
  wire       [0:0]    stage0_dataColisions;
  wire       [0:0]    stage0_wayInvalidate;
  wire                stage0_isAmo;
  wire                when_DataCache_l771;
  reg                 stageA_request_wr;
  reg        [1:0]    stageA_request_size;
  reg                 stageA_request_totalyConsistent;
  wire                when_DataCache_l771_1;
  reg        [3:0]    stageA_mask;
  wire                stageA_isAmo;
  wire                stageA_isLrsc;
  wire       [0:0]    stageA_wayHits;
  wire                when_DataCache_l771_2;
  reg        [0:0]    stageA_wayInvalidate;
  wire                when_DataCache_l771_3;
  reg        [0:0]    stage0_dataColisions_regNextWhen;
  wire       [0:0]    _zz_stageA_dataColisions;
  wire       [0:0]    stageA_dataColisions;
  wire                when_DataCache_l822;
  reg                 stageB_request_wr;
  reg        [1:0]    stageB_request_size;
  reg                 stageB_request_totalyConsistent;
  reg                 stageB_mmuRspFreeze;
  wire                when_DataCache_l824;
  reg        [31:0]   stageB_mmuRsp_physicalAddress;
  reg                 stageB_mmuRsp_isIoAccess;
  reg                 stageB_mmuRsp_isPaging;
  reg                 stageB_mmuRsp_allowRead;
  reg                 stageB_mmuRsp_allowWrite;
  reg                 stageB_mmuRsp_allowExecute;
  reg                 stageB_mmuRsp_exception;
  reg                 stageB_mmuRsp_refilling;
  reg                 stageB_mmuRsp_bypassTranslation;
  wire                when_DataCache_l821;
  reg                 stageB_tagsReadRsp_0_valid;
  reg                 stageB_tagsReadRsp_0_error;
  reg        [19:0]   stageB_tagsReadRsp_0_address;
  wire                when_DataCache_l821_1;
  reg        [31:0]   stageB_dataReadRsp_0;
  wire                when_DataCache_l820;
  reg        [0:0]    stageB_wayInvalidate;
  wire                stageB_consistancyHazard;
  wire                when_DataCache_l820_1;
  reg        [0:0]    stageB_dataColisions;
  wire                when_DataCache_l820_2;
  reg                 stageB_unaligned;
  wire                when_DataCache_l820_3;
  reg        [0:0]    stageB_waysHitsBeforeInvalidate;
  wire       [0:0]    stageB_waysHits;
  wire                stageB_waysHit;
  wire       [31:0]   stageB_dataMux;
  wire                when_DataCache_l820_4;
  reg        [3:0]    stageB_mask;
  reg                 stageB_loaderValid;
  wire       [31:0]   stageB_ioMemRspMuxed;
  reg                 stageB_flusher_waitDone;
  wire                stageB_flusher_hold;
  reg        [7:0]    stageB_flusher_counter;
  wire                when_DataCache_l850;
  wire                when_DataCache_l856;
  reg                 stageB_flusher_start;
  wire                stageB_isAmo;
  wire                stageB_isAmoCached;
  wire                stageB_isExternalLsrc;
  wire                stageB_isExternalAmo;
  wire       [31:0]   stageB_requestDataBypass;
  reg                 stageB_cpuWriteToCache;
  wire                when_DataCache_l926;
  wire                stageB_badPermissions;
  wire                stageB_loadStoreFault;
  wire                stageB_bypassCache;
  wire                when_DataCache_l995;
  wire                when_DataCache_l1004;
  wire                when_DataCache_l1009;
  wire                when_DataCache_l1020;
  wire                when_DataCache_l1032;
  wire                when_DataCache_l991;
  wire                when_DataCache_l1066;
  wire                when_DataCache_l1075;
  reg                 loader_valid;
  reg                 loader_counter_willIncrement;
  wire                loader_counter_willClear;
  reg        [2:0]    loader_counter_valueNext;
  reg        [2:0]    loader_counter_value;
  wire                loader_counter_willOverflowIfInc;
  wire                loader_counter_willOverflow;
  reg        [0:0]    loader_waysAllocator;
  reg                 loader_error;
  wire                loader_kill;
  reg                 loader_killReg;
  wire                when_DataCache_l1090;
  wire                loader_done;
  wire                when_DataCache_l1118;
  reg                 loader_valid_regNext;
  wire                when_DataCache_l1122;
  wire                when_DataCache_l1125;
  (* no_rw_check , ram_style = "block" *) reg [21:0] ways_0_tags [0:127];
  (* no_rw_check , ram_style = "block" *) reg [7:0] ways_0_data_symbol0 [0:1023];
  (* no_rw_check , ram_style = "block" *) reg [7:0] ways_0_data_symbol1 [0:1023];
  (* no_rw_check , ram_style = "block" *) reg [7:0] ways_0_data_symbol2 [0:1023];
  (* no_rw_check , ram_style = "block" *) reg [7:0] ways_0_data_symbol3 [0:1023];
  reg [7:0] _zz_ways_0_datasymbol_read;
  reg [7:0] _zz_ways_0_datasymbol_read_1;
  reg [7:0] _zz_ways_0_datasymbol_read_2;
  reg [7:0] _zz_ways_0_datasymbol_read_3;

  assign _zz_stage0_dataColisions = (io_cpu_execute_address[11 : 2] >>> 0);
  assign _zz__zz_stageA_dataColisions = (io_cpu_memory_address[11 : 2] >>> 0);
  assign _zz_when = 1'b1;
  assign _zz_loader_counter_valueNext_1 = loader_counter_willIncrement;
  assign _zz_loader_counter_valueNext = {2'd0, _zz_loader_counter_valueNext_1};
  assign _zz_loader_waysAllocator = {loader_waysAllocator,loader_waysAllocator[0]};
  assign _zz_ways_0_tags_port = {tagsWriteCmd_payload_data_address,{tagsWriteCmd_payload_data_error,tagsWriteCmd_payload_data_valid}};
  always @(posedge clk) begin
    if(_zz_ways_0_tagsReadRsp_valid) begin
      _zz_ways_0_tags_port0 <= ways_0_tags[tagsReadCmd_payload];
    end
  end

  always @(posedge clk) begin
    if(_zz_2) begin
      ways_0_tags[tagsWriteCmd_payload_address] <= _zz_ways_0_tags_port;
    end
  end

  always @(*) begin
    _zz_ways_0_data_port0 = {_zz_ways_0_datasymbol_read_3, _zz_ways_0_datasymbol_read_2, _zz_ways_0_datasymbol_read_1, _zz_ways_0_datasymbol_read};
  end
  always @(posedge clk) begin
    if(_zz_ways_0_dataReadRspMem) begin
      _zz_ways_0_datasymbol_read <= ways_0_data_symbol0[dataReadCmd_payload];
      _zz_ways_0_datasymbol_read_1 <= ways_0_data_symbol1[dataReadCmd_payload];
      _zz_ways_0_datasymbol_read_2 <= ways_0_data_symbol2[dataReadCmd_payload];
      _zz_ways_0_datasymbol_read_3 <= ways_0_data_symbol3[dataReadCmd_payload];
    end
  end

  always @(posedge clk) begin
    if(dataWriteCmd_payload_mask[0] && _zz_1) begin
      ways_0_data_symbol0[dataWriteCmd_payload_address] <= dataWriteCmd_payload_data[7 : 0];
    end
    if(dataWriteCmd_payload_mask[1] && _zz_1) begin
      ways_0_data_symbol1[dataWriteCmd_payload_address] <= dataWriteCmd_payload_data[15 : 8];
    end
    if(dataWriteCmd_payload_mask[2] && _zz_1) begin
      ways_0_data_symbol2[dataWriteCmd_payload_address] <= dataWriteCmd_payload_data[23 : 16];
    end
    if(dataWriteCmd_payload_mask[3] && _zz_1) begin
      ways_0_data_symbol3[dataWriteCmd_payload_address] <= dataWriteCmd_payload_data[31 : 24];
    end
  end

  always @(*) begin
    _zz_1 = 1'b0;
    if(when_DataCache_l645) begin
      _zz_1 = 1'b1;
    end
  end

  always @(*) begin
    _zz_2 = 1'b0;
    if(when_DataCache_l642) begin
      _zz_2 = 1'b1;
    end
  end

  assign haltCpu = 1'b0;
  assign _zz_ways_0_tagsReadRsp_valid = (tagsReadCmd_valid && (! io_cpu_memory_isStuck));
  assign _zz_ways_0_tagsReadRsp_valid_1 = _zz_ways_0_tags_port0;
  assign ways_0_tagsReadRsp_valid = _zz_ways_0_tagsReadRsp_valid_1[0];
  assign ways_0_tagsReadRsp_error = _zz_ways_0_tagsReadRsp_valid_1[1];
  assign ways_0_tagsReadRsp_address = _zz_ways_0_tagsReadRsp_valid_1[21 : 2];
  assign _zz_ways_0_dataReadRspMem = (dataReadCmd_valid && (! io_cpu_memory_isStuck));
  assign ways_0_dataReadRspMem = _zz_ways_0_data_port0;
  assign ways_0_dataReadRsp = ways_0_dataReadRspMem[31 : 0];
  assign when_DataCache_l642 = (tagsWriteCmd_valid && tagsWriteCmd_payload_way[0]);
  assign when_DataCache_l645 = (dataWriteCmd_valid && dataWriteCmd_payload_way[0]);
  always @(*) begin
    tagsReadCmd_valid = 1'b0;
    if(when_DataCache_l664) begin
      tagsReadCmd_valid = 1'b1;
    end
  end

  always @(*) begin
    tagsReadCmd_payload = 7'bxxxxxxx;
    if(when_DataCache_l664) begin
      tagsReadCmd_payload = io_cpu_execute_address[11 : 5];
    end
  end

  always @(*) begin
    dataReadCmd_valid = 1'b0;
    if(when_DataCache_l664) begin
      dataReadCmd_valid = 1'b1;
    end
  end

  always @(*) begin
    dataReadCmd_payload = 10'bxxxxxxxxxx;
    if(when_DataCache_l664) begin
      dataReadCmd_payload = io_cpu_execute_address[11 : 2];
    end
  end

  always @(*) begin
    tagsWriteCmd_valid = 1'b0;
    if(when_DataCache_l850) begin
      tagsWriteCmd_valid = 1'b1;
    end
    if(when_DataCache_l1066) begin
      tagsWriteCmd_valid = 1'b0;
    end
    if(loader_done) begin
      tagsWriteCmd_valid = 1'b1;
    end
  end

  always @(*) begin
    tagsWriteCmd_payload_way = 1'bx;
    if(when_DataCache_l850) begin
      tagsWriteCmd_payload_way = 1'b1;
    end
    if(loader_done) begin
      tagsWriteCmd_payload_way = loader_waysAllocator;
    end
  end

  always @(*) begin
    tagsWriteCmd_payload_address = 7'bxxxxxxx;
    if(when_DataCache_l850) begin
      tagsWriteCmd_payload_address = stageB_flusher_counter[6:0];
    end
    if(loader_done) begin
      tagsWriteCmd_payload_address = stageB_mmuRsp_physicalAddress[11 : 5];
    end
  end

  always @(*) begin
    tagsWriteCmd_payload_data_valid = 1'bx;
    if(when_DataCache_l850) begin
      tagsWriteCmd_payload_data_valid = 1'b0;
    end
    if(loader_done) begin
      tagsWriteCmd_payload_data_valid = (! (loader_kill || loader_killReg));
    end
  end

  always @(*) begin
    tagsWriteCmd_payload_data_error = 1'bx;
    if(loader_done) begin
      tagsWriteCmd_payload_data_error = (loader_error || (io_mem_rsp_valid && io_mem_rsp_payload_error));
    end
  end

  always @(*) begin
    tagsWriteCmd_payload_data_address = 20'bxxxxxxxxxxxxxxxxxxxx;
    if(loader_done) begin
      tagsWriteCmd_payload_data_address = stageB_mmuRsp_physicalAddress[31 : 12];
    end
  end

  always @(*) begin
    dataWriteCmd_valid = 1'b0;
    if(stageB_cpuWriteToCache) begin
      if(when_DataCache_l926) begin
        dataWriteCmd_valid = 1'b1;
      end
    end
    if(when_DataCache_l1066) begin
      dataWriteCmd_valid = 1'b0;
    end
    if(when_DataCache_l1090) begin
      dataWriteCmd_valid = 1'b1;
    end
  end

  always @(*) begin
    dataWriteCmd_payload_way = 1'bx;
    if(stageB_cpuWriteToCache) begin
      dataWriteCmd_payload_way = stageB_waysHits;
    end
    if(when_DataCache_l1090) begin
      dataWriteCmd_payload_way = loader_waysAllocator;
    end
  end

  always @(*) begin
    dataWriteCmd_payload_address = 10'bxxxxxxxxxx;
    if(stageB_cpuWriteToCache) begin
      dataWriteCmd_payload_address = stageB_mmuRsp_physicalAddress[11 : 2];
    end
    if(when_DataCache_l1090) begin
      dataWriteCmd_payload_address = {stageB_mmuRsp_physicalAddress[11 : 5],loader_counter_value};
    end
  end

  always @(*) begin
    dataWriteCmd_payload_data = 32'bxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxxx;
    if(stageB_cpuWriteToCache) begin
      dataWriteCmd_payload_data[31 : 0] = stageB_requestDataBypass;
    end
    if(when_DataCache_l1090) begin
      dataWriteCmd_payload_data = io_mem_rsp_payload_data;
    end
  end

  always @(*) begin
    dataWriteCmd_payload_mask = 4'bxxxx;
    if(stageB_cpuWriteToCache) begin
      dataWriteCmd_payload_mask = 4'b0000;
      if(_zz_when[0]) begin
        dataWriteCmd_payload_mask[3 : 0] = stageB_mask;
      end
    end
    if(when_DataCache_l1090) begin
      dataWriteCmd_payload_mask = 4'b1111;
    end
  end

  assign when_DataCache_l664 = (io_cpu_execute_isValid && (! io_cpu_memory_isStuck));
  always @(*) begin
    io_cpu_execute_haltIt = 1'b0;
    if(when_DataCache_l850) begin
      io_cpu_execute_haltIt = 1'b1;
    end
  end

  assign rspSync = 1'b1;
  assign rspLast = 1'b1;
  assign io_mem_cmd_fire = (io_mem_cmd_valid && io_mem_cmd_ready);
  assign when_DataCache_l686 = (! io_cpu_writeBack_isStuck);
  always @(*) begin
    _zz_stage0_mask = 4'bxxxx;
    case(io_cpu_execute_args_size)
      2'b00 : begin
        _zz_stage0_mask = 4'b0001;
      end
      2'b01 : begin
        _zz_stage0_mask = 4'b0011;
      end
      2'b10 : begin
        _zz_stage0_mask = 4'b1111;
      end
      default : begin
      end
    endcase
  end

  assign stage0_mask = (_zz_stage0_mask <<< io_cpu_execute_address[1 : 0]);
  assign stage0_dataColisions[0] = (((dataWriteCmd_valid && dataWriteCmd_payload_way[0]) && (dataWriteCmd_payload_address == _zz_stage0_dataColisions)) && ((stage0_mask & dataWriteCmd_payload_mask[3 : 0]) != 4'b0000));
  assign stage0_wayInvalidate = 1'b0;
  assign stage0_isAmo = 1'b0;
  assign when_DataCache_l771 = (! io_cpu_memory_isStuck);
  assign when_DataCache_l771_1 = (! io_cpu_memory_isStuck);
  assign io_cpu_memory_isWrite = stageA_request_wr;
  assign stageA_isAmo = 1'b0;
  assign stageA_isLrsc = 1'b0;
  assign stageA_wayHits = ((io_cpu_memory_mmuRsp_physicalAddress[31 : 12] == ways_0_tagsReadRsp_address) && ways_0_tagsReadRsp_valid);
  assign when_DataCache_l771_2 = (! io_cpu_memory_isStuck);
  assign when_DataCache_l771_3 = (! io_cpu_memory_isStuck);
  assign _zz_stageA_dataColisions[0] = (((dataWriteCmd_valid && dataWriteCmd_payload_way[0]) && (dataWriteCmd_payload_address == _zz__zz_stageA_dataColisions)) && ((stageA_mask & dataWriteCmd_payload_mask[3 : 0]) != 4'b0000));
  assign stageA_dataColisions = (stage0_dataColisions_regNextWhen | _zz_stageA_dataColisions);
  assign when_DataCache_l822 = (! io_cpu_writeBack_isStuck);
  always @(*) begin
    stageB_mmuRspFreeze = 1'b0;
    if(when_DataCache_l1125) begin
      stageB_mmuRspFreeze = 1'b1;
    end
  end

  assign when_DataCache_l824 = ((! io_cpu_writeBack_isStuck) && (! stageB_mmuRspFreeze));
  assign when_DataCache_l821 = (! io_cpu_writeBack_isStuck);
  assign when_DataCache_l821_1 = (! io_cpu_writeBack_isStuck);
  assign when_DataCache_l820 = (! io_cpu_writeBack_isStuck);
  assign stageB_consistancyHazard = 1'b0;
  assign when_DataCache_l820_1 = (! io_cpu_writeBack_isStuck);
  assign when_DataCache_l820_2 = (! io_cpu_writeBack_isStuck);
  assign when_DataCache_l820_3 = (! io_cpu_writeBack_isStuck);
  assign stageB_waysHits = (stageB_waysHitsBeforeInvalidate & (~ stageB_wayInvalidate));
  assign stageB_waysHit = (|stageB_waysHits);
  assign stageB_dataMux = stageB_dataReadRsp_0;
  assign when_DataCache_l820_4 = (! io_cpu_writeBack_isStuck);
  always @(*) begin
    stageB_loaderValid = 1'b0;
    if(io_cpu_writeBack_isValid) begin
      if(!stageB_isExternalAmo) begin
        if(!when_DataCache_l991) begin
          if(!when_DataCache_l1004) begin
            if(io_mem_cmd_ready) begin
              stageB_loaderValid = 1'b1;
            end
          end
        end
      end
    end
    if(when_DataCache_l1066) begin
      stageB_loaderValid = 1'b0;
    end
  end

  assign stageB_ioMemRspMuxed = io_mem_rsp_payload_data[31 : 0];
  always @(*) begin
    io_cpu_writeBack_haltIt = 1'b1;
    if(io_cpu_writeBack_isValid) begin
      if(!stageB_isExternalAmo) begin
        if(when_DataCache_l991) begin
          if(when_DataCache_l995) begin
            io_cpu_writeBack_haltIt = 1'b0;
          end
        end else begin
          if(when_DataCache_l1004) begin
            if(when_DataCache_l1009) begin
              io_cpu_writeBack_haltIt = 1'b0;
            end
          end
        end
      end
    end
    if(when_DataCache_l1066) begin
      io_cpu_writeBack_haltIt = 1'b0;
    end
  end

  assign stageB_flusher_hold = 1'b0;
  assign when_DataCache_l850 = (! stageB_flusher_counter[7]);
  assign when_DataCache_l856 = (! stageB_flusher_hold);
  assign io_cpu_flush_ready = (stageB_flusher_waitDone && stageB_flusher_counter[7]);
  assign stageB_isAmo = 1'b0;
  assign stageB_isAmoCached = 1'b0;
  assign stageB_isExternalLsrc = 1'b0;
  assign stageB_isExternalAmo = 1'b0;
  assign stageB_requestDataBypass = io_cpu_writeBack_storeData;
  always @(*) begin
    stageB_cpuWriteToCache = 1'b0;
    if(io_cpu_writeBack_isValid) begin
      if(!stageB_isExternalAmo) begin
        if(!when_DataCache_l991) begin
          if(when_DataCache_l1004) begin
            stageB_cpuWriteToCache = 1'b1;
          end
        end
      end
    end
  end

  assign when_DataCache_l926 = (stageB_request_wr && stageB_waysHit);
  assign stageB_badPermissions = (((! stageB_mmuRsp_allowWrite) && stageB_request_wr) || ((! stageB_mmuRsp_allowRead) && ((! stageB_request_wr) || stageB_isAmo)));
  assign stageB_loadStoreFault = (io_cpu_writeBack_isValid && (stageB_mmuRsp_exception || stageB_badPermissions));
  always @(*) begin
    io_cpu_redo = 1'b0;
    if(io_cpu_writeBack_isValid) begin
      if(!stageB_isExternalAmo) begin
        if(!when_DataCache_l991) begin
          if(when_DataCache_l1004) begin
            if(when_DataCache_l1020) begin
              io_cpu_redo = 1'b1;
            end
          end
        end
      end
    end
    if(when_DataCache_l1075) begin
      io_cpu_redo = 1'b1;
    end
    if(when_DataCache_l1122) begin
      io_cpu_redo = 1'b1;
    end
  end

  always @(*) begin
    io_cpu_writeBack_accessError = 1'b0;
    if(stageB_bypassCache) begin
      io_cpu_writeBack_accessError = ((((! stageB_request_wr) && 1'b1) && io_mem_rsp_valid) && io_mem_rsp_payload_error);
    end else begin
      io_cpu_writeBack_accessError = (((stageB_waysHits & stageB_tagsReadRsp_0_error) != 1'b0) || (stageB_loadStoreFault && (! stageB_mmuRsp_isPaging)));
    end
  end

  assign io_cpu_writeBack_mmuException = (stageB_loadStoreFault && stageB_mmuRsp_isPaging);
  assign io_cpu_writeBack_unalignedAccess = (io_cpu_writeBack_isValid && stageB_unaligned);
  assign io_cpu_writeBack_isWrite = stageB_request_wr;
  always @(*) begin
    io_mem_cmd_valid = 1'b0;
    if(io_cpu_writeBack_isValid) begin
      if(!stageB_isExternalAmo) begin
        if(when_DataCache_l991) begin
          io_mem_cmd_valid = (! memCmdSent);
        end else begin
          if(when_DataCache_l1004) begin
            if(stageB_request_wr) begin
              io_mem_cmd_valid = 1'b1;
            end
          end else begin
            if(when_DataCache_l1032) begin
              io_mem_cmd_valid = 1'b1;
            end
          end
        end
      end
    end
    if(when_DataCache_l1066) begin
      io_mem_cmd_valid = 1'b0;
    end
  end

  always @(*) begin
    io_mem_cmd_payload_address = stageB_mmuRsp_physicalAddress;
    if(io_cpu_writeBack_isValid) begin
      if(!stageB_isExternalAmo) begin
        if(!when_DataCache_l991) begin
          if(!when_DataCache_l1004) begin
            io_mem_cmd_payload_address[4 : 0] = 5'h0;
          end
        end
      end
    end
  end

  assign io_mem_cmd_payload_last = 1'b1;
  always @(*) begin
    io_mem_cmd_payload_wr = stageB_request_wr;
    if(io_cpu_writeBack_isValid) begin
      if(!stageB_isExternalAmo) begin
        if(!when_DataCache_l991) begin
          if(!when_DataCache_l1004) begin
            io_mem_cmd_payload_wr = 1'b0;
          end
        end
      end
    end
  end

  assign io_mem_cmd_payload_mask = stageB_mask;
  assign io_mem_cmd_payload_data = stageB_requestDataBypass;
  assign io_mem_cmd_payload_uncached = stageB_mmuRsp_isIoAccess;
  always @(*) begin
    io_mem_cmd_payload_size = {1'd0, stageB_request_size};
    if(io_cpu_writeBack_isValid) begin
      if(!stageB_isExternalAmo) begin
        if(!when_DataCache_l991) begin
          if(!when_DataCache_l1004) begin
            io_mem_cmd_payload_size = 3'b101;
          end
        end
      end
    end
  end

  assign stageB_bypassCache = ((stageB_mmuRsp_isIoAccess || stageB_isExternalLsrc) || stageB_isExternalAmo);
  assign io_cpu_writeBack_keepMemRspData = 1'b0;
  assign when_DataCache_l995 = ((! stageB_request_wr) ? (io_mem_rsp_valid && rspSync) : io_mem_cmd_ready);
  assign when_DataCache_l1004 = (stageB_waysHit || (stageB_request_wr && (! stageB_isAmoCached)));
  assign when_DataCache_l1009 = ((! stageB_request_wr) || io_mem_cmd_ready);
  assign when_DataCache_l1020 = (((! stageB_request_wr) || stageB_isAmoCached) && ((stageB_dataColisions & stageB_waysHits) != 1'b0));
  assign when_DataCache_l1032 = (! memCmdSent);
  assign when_DataCache_l991 = (stageB_mmuRsp_isIoAccess || stageB_isExternalLsrc);
  always @(*) begin
    if(stageB_bypassCache) begin
      io_cpu_writeBack_data = stageB_ioMemRspMuxed;
    end else begin
      io_cpu_writeBack_data = stageB_dataMux;
    end
  end

  assign when_DataCache_l1066 = ((((stageB_consistancyHazard || stageB_mmuRsp_refilling) || io_cpu_writeBack_accessError) || io_cpu_writeBack_mmuException) || io_cpu_writeBack_unalignedAccess);
  assign when_DataCache_l1075 = (io_cpu_writeBack_isValid && (stageB_mmuRsp_refilling || stageB_consistancyHazard));
  always @(*) begin
    loader_counter_willIncrement = 1'b0;
    if(when_DataCache_l1090) begin
      loader_counter_willIncrement = 1'b1;
    end
  end

  assign loader_counter_willClear = 1'b0;
  assign loader_counter_willOverflowIfInc = (loader_counter_value == 3'b111);
  assign loader_counter_willOverflow = (loader_counter_willOverflowIfInc && loader_counter_willIncrement);
  always @(*) begin
    loader_counter_valueNext = (loader_counter_value + _zz_loader_counter_valueNext);
    if(loader_counter_willClear) begin
      loader_counter_valueNext = 3'b000;
    end
  end

  assign loader_kill = 1'b0;
  assign when_DataCache_l1090 = ((loader_valid && io_mem_rsp_valid) && rspLast);
  assign loader_done = loader_counter_willOverflow;
  assign when_DataCache_l1118 = (! loader_valid);
  assign when_DataCache_l1122 = (loader_valid && (! loader_valid_regNext));
  assign io_cpu_execute_refilling = loader_valid;
  assign when_DataCache_l1125 = (stageB_loaderValid || loader_valid);
  always @(posedge clk) begin
    tagsWriteLastCmd_valid <= tagsWriteCmd_valid;
    tagsWriteLastCmd_payload_way <= tagsWriteCmd_payload_way;
    tagsWriteLastCmd_payload_address <= tagsWriteCmd_payload_address;
    tagsWriteLastCmd_payload_data_valid <= tagsWriteCmd_payload_data_valid;
    tagsWriteLastCmd_payload_data_error <= tagsWriteCmd_payload_data_error;
    tagsWriteLastCmd_payload_data_address <= tagsWriteCmd_payload_data_address;
    if(when_DataCache_l771) begin
      stageA_request_wr <= io_cpu_execute_args_wr;
      stageA_request_size <= io_cpu_execute_args_size;
      stageA_request_totalyConsistent <= io_cpu_execute_args_totalyConsistent;
    end
    if(when_DataCache_l771_1) begin
      stageA_mask <= stage0_mask;
    end
    if(when_DataCache_l771_2) begin
      stageA_wayInvalidate <= stage0_wayInvalidate;
    end
    if(when_DataCache_l771_3) begin
      stage0_dataColisions_regNextWhen <= stage0_dataColisions;
    end
    if(when_DataCache_l822) begin
      stageB_request_wr <= stageA_request_wr;
      stageB_request_size <= stageA_request_size;
      stageB_request_totalyConsistent <= stageA_request_totalyConsistent;
    end
    if(when_DataCache_l824) begin
      stageB_mmuRsp_physicalAddress <= io_cpu_memory_mmuRsp_physicalAddress;
      stageB_mmuRsp_isIoAccess <= io_cpu_memory_mmuRsp_isIoAccess;
      stageB_mmuRsp_isPaging <= io_cpu_memory_mmuRsp_isPaging;
      stageB_mmuRsp_allowRead <= io_cpu_memory_mmuRsp_allowRead;
      stageB_mmuRsp_allowWrite <= io_cpu_memory_mmuRsp_allowWrite;
      stageB_mmuRsp_allowExecute <= io_cpu_memory_mmuRsp_allowExecute;
      stageB_mmuRsp_exception <= io_cpu_memory_mmuRsp_exception;
      stageB_mmuRsp_refilling <= io_cpu_memory_mmuRsp_refilling;
      stageB_mmuRsp_bypassTranslation <= io_cpu_memory_mmuRsp_bypassTranslation;
    end
    if(when_DataCache_l821) begin
      stageB_tagsReadRsp_0_valid <= ways_0_tagsReadRsp_valid;
      stageB_tagsReadRsp_0_error <= ways_0_tagsReadRsp_error;
      stageB_tagsReadRsp_0_address <= ways_0_tagsReadRsp_address;
    end
    if(when_DataCache_l821_1) begin
      stageB_dataReadRsp_0 <= ways_0_dataReadRsp;
    end
    if(when_DataCache_l820) begin
      stageB_wayInvalidate <= stageA_wayInvalidate;
    end
    if(when_DataCache_l820_1) begin
      stageB_dataColisions <= stageA_dataColisions;
    end
    if(when_DataCache_l820_2) begin
      stageB_unaligned <= ({((stageA_request_size == 2'b10) && (io_cpu_memory_address[1 : 0] != 2'b00)),((stageA_request_size == 2'b01) && (io_cpu_memory_address[0 : 0] != 1'b0))} != 2'b00);
    end
    if(when_DataCache_l820_3) begin
      stageB_waysHitsBeforeInvalidate <= stageA_wayHits;
    end
    if(when_DataCache_l820_4) begin
      stageB_mask <= stageA_mask;
    end
    loader_valid_regNext <= loader_valid;
  end

  always @(posedge clk) begin
    if(reset) begin
      memCmdSent <= 1'b0;
      stageB_flusher_waitDone <= 1'b0;
      stageB_flusher_counter <= 8'h0;
      stageB_flusher_start <= 1'b1;
      loader_valid <= 1'b0;
      loader_counter_value <= 3'b000;
      loader_waysAllocator <= 1'b1;
      loader_error <= 1'b0;
      loader_killReg <= 1'b0;
    end else begin
      if(io_mem_cmd_fire) begin
        memCmdSent <= 1'b1;
      end
      if(when_DataCache_l686) begin
        memCmdSent <= 1'b0;
      end
      if(io_cpu_flush_ready) begin
        stageB_flusher_waitDone <= 1'b0;
      end
      if(when_DataCache_l850) begin
        if(when_DataCache_l856) begin
          stageB_flusher_counter <= (stageB_flusher_counter + 8'h01);
          if(io_cpu_flush_payload_singleLine) begin
            stageB_flusher_counter[7] <= 1'b1;
          end
        end
      end
      stageB_flusher_start <= (((((((! stageB_flusher_waitDone) && (! stageB_flusher_start)) && io_cpu_flush_valid) && (! io_cpu_execute_isValid)) && (! io_cpu_memory_isValid)) && (! io_cpu_writeBack_isValid)) && (! io_cpu_redo));
      if(stageB_flusher_start) begin
        stageB_flusher_waitDone <= 1'b1;
        stageB_flusher_counter <= 8'h0;
        if(io_cpu_flush_payload_singleLine) begin
          stageB_flusher_counter <= {1'b0,io_cpu_flush_payload_lineId};
        end
      end
      `ifndef SYNTHESIS
        `ifdef FORMAL
          assert((! ((io_cpu_writeBack_isValid && (! io_cpu_writeBack_haltIt)) && io_cpu_writeBack_isStuck))); // DataCache.scala:L1077
        `else
          if(!(! ((io_cpu_writeBack_isValid && (! io_cpu_writeBack_haltIt)) && io_cpu_writeBack_isStuck))) begin
            $display("ERROR writeBack stuck by another plugin is not allowed"); // DataCache.scala:L1077
          end
        `endif
      `endif
      if(stageB_loaderValid) begin
        loader_valid <= 1'b1;
      end
      loader_counter_value <= loader_counter_valueNext;
      if(loader_kill) begin
        loader_killReg <= 1'b1;
      end
      if(when_DataCache_l1090) begin
        loader_error <= (loader_error || io_mem_rsp_payload_error);
      end
      if(loader_done) begin
        loader_valid <= 1'b0;
        loader_error <= 1'b0;
        loader_killReg <= 1'b0;
      end
      if(when_DataCache_l1118) begin
        loader_waysAllocator <= _zz_loader_waysAllocator[0:0];
      end
    end
  end


endmodule

module InstructionCache (
  input               io_flush,
  input               io_cpu_prefetch_isValid,
  output reg          io_cpu_prefetch_haltIt,
  input      [31:0]   io_cpu_prefetch_pc,
  input               io_cpu_fetch_isValid,
  input               io_cpu_fetch_isStuck,
  input               io_cpu_fetch_isRemoved,
  input      [31:0]   io_cpu_fetch_pc,
  output     [31:0]   io_cpu_fetch_data,
  input      [31:0]   io_cpu_fetch_mmuRsp_physicalAddress,
  input               io_cpu_fetch_mmuRsp_isIoAccess,
  input               io_cpu_fetch_mmuRsp_isPaging,
  input               io_cpu_fetch_mmuRsp_allowRead,
  input               io_cpu_fetch_mmuRsp_allowWrite,
  input               io_cpu_fetch_mmuRsp_allowExecute,
  input               io_cpu_fetch_mmuRsp_exception,
  input               io_cpu_fetch_mmuRsp_refilling,
  input               io_cpu_fetch_mmuRsp_bypassTranslation,
  output     [31:0]   io_cpu_fetch_physicalAddress,
  input               io_cpu_decode_isValid,
  input               io_cpu_decode_isStuck,
  input      [31:0]   io_cpu_decode_pc,
  output     [31:0]   io_cpu_decode_physicalAddress,
  output     [31:0]   io_cpu_decode_data,
  output              io_cpu_decode_cacheMiss,
  output              io_cpu_decode_error,
  output              io_cpu_decode_mmuRefilling,
  output              io_cpu_decode_mmuException,
  input               io_cpu_decode_isUser,
  input               io_cpu_fill_valid,
  input      [31:0]   io_cpu_fill_payload,
  output              io_mem_cmd_valid,
  input               io_mem_cmd_ready,
  output     [31:0]   io_mem_cmd_payload_address,
  output     [2:0]    io_mem_cmd_payload_size,
  input               io_mem_rsp_valid,
  input      [31:0]   io_mem_rsp_payload_data,
  input               io_mem_rsp_payload_error,
  input               clk,
  input               reset
);

  reg        [31:0]   _zz_banks_0_port1;
  reg        [21:0]   _zz_ways_0_tags_port1;
  wire       [21:0]   _zz_ways_0_tags_port;
  reg                 _zz_1;
  reg                 _zz_2;
  reg                 lineLoader_fire;
  reg                 lineLoader_valid;
  (* keep , syn_keep *) reg        [31:0]   lineLoader_address /* synthesis syn_keep = 1 */ ;
  reg                 lineLoader_hadError;
  reg                 lineLoader_flushPending;
  reg        [7:0]    lineLoader_flushCounter;
  wire                when_InstructionCache_l338;
  reg                 _zz_when_InstructionCache_l342;
  wire                when_InstructionCache_l342;
  wire                when_InstructionCache_l351;
  reg                 lineLoader_cmdSent;
  wire                io_mem_cmd_fire;
  wire                when_Utils_l515;
  reg                 lineLoader_wayToAllocate_willIncrement;
  wire                lineLoader_wayToAllocate_willClear;
  wire                lineLoader_wayToAllocate_willOverflowIfInc;
  wire                lineLoader_wayToAllocate_willOverflow;
  (* keep , syn_keep *) reg        [2:0]    lineLoader_wordIndex /* synthesis syn_keep = 1 */ ;
  wire                lineLoader_write_tag_0_valid;
  wire       [6:0]    lineLoader_write_tag_0_payload_address;
  wire                lineLoader_write_tag_0_payload_data_valid;
  wire                lineLoader_write_tag_0_payload_data_error;
  wire       [19:0]   lineLoader_write_tag_0_payload_data_address;
  wire                lineLoader_write_data_0_valid;
  wire       [9:0]    lineLoader_write_data_0_payload_address;
  wire       [31:0]   lineLoader_write_data_0_payload_data;
  wire                when_InstructionCache_l401;
  wire       [9:0]    _zz_fetchStage_read_banksValue_0_dataMem;
  wire                _zz_fetchStage_read_banksValue_0_dataMem_1;
  wire       [31:0]   fetchStage_read_banksValue_0_dataMem;
  wire       [31:0]   fetchStage_read_banksValue_0_data;
  wire       [6:0]    _zz_fetchStage_read_waysValues_0_tag_valid;
  wire                _zz_fetchStage_read_waysValues_0_tag_valid_1;
  wire                fetchStage_read_waysValues_0_tag_valid;
  wire                fetchStage_read_waysValues_0_tag_error;
  wire       [19:0]   fetchStage_read_waysValues_0_tag_address;
  wire       [21:0]   _zz_fetchStage_read_waysValues_0_tag_valid_2;
  wire                fetchStage_hit_hits_0;
  wire                fetchStage_hit_valid;
  wire                fetchStage_hit_error;
  wire       [31:0]   fetchStage_hit_data;
  wire       [31:0]   fetchStage_hit_word;
  wire                when_InstructionCache_l435;
  reg        [31:0]   io_cpu_fetch_data_regNextWhen;
  wire                when_InstructionCache_l459;
  reg        [31:0]   decodeStage_mmuRsp_physicalAddress;
  reg                 decodeStage_mmuRsp_isIoAccess;
  reg                 decodeStage_mmuRsp_isPaging;
  reg                 decodeStage_mmuRsp_allowRead;
  reg                 decodeStage_mmuRsp_allowWrite;
  reg                 decodeStage_mmuRsp_allowExecute;
  reg                 decodeStage_mmuRsp_exception;
  reg                 decodeStage_mmuRsp_refilling;
  reg                 decodeStage_mmuRsp_bypassTranslation;
  wire                when_InstructionCache_l459_1;
  reg                 decodeStage_hit_valid;
  wire                when_InstructionCache_l459_2;
  reg                 decodeStage_hit_error;
  (* no_rw_check , ram_style = "block" *) reg [31:0] banks_0 [0:1023];
  (* no_rw_check , ram_style = "block" *) reg [21:0] ways_0_tags [0:127];

  assign _zz_ways_0_tags_port = {lineLoader_write_tag_0_payload_data_address,{lineLoader_write_tag_0_payload_data_error,lineLoader_write_tag_0_payload_data_valid}};
  always @(posedge clk) begin
    if(_zz_1) begin
      banks_0[lineLoader_write_data_0_payload_address] <= lineLoader_write_data_0_payload_data;
    end
  end

  always @(posedge clk) begin
    if(_zz_fetchStage_read_banksValue_0_dataMem_1) begin
      _zz_banks_0_port1 <= banks_0[_zz_fetchStage_read_banksValue_0_dataMem];
    end
  end

  always @(posedge clk) begin
    if(_zz_2) begin
      ways_0_tags[lineLoader_write_tag_0_payload_address] <= _zz_ways_0_tags_port;
    end
  end

  always @(posedge clk) begin
    if(_zz_fetchStage_read_waysValues_0_tag_valid_1) begin
      _zz_ways_0_tags_port1 <= ways_0_tags[_zz_fetchStage_read_waysValues_0_tag_valid];
    end
  end

  always @(*) begin
    _zz_1 = 1'b0;
    if(lineLoader_write_data_0_valid) begin
      _zz_1 = 1'b1;
    end
  end

  always @(*) begin
    _zz_2 = 1'b0;
    if(lineLoader_write_tag_0_valid) begin
      _zz_2 = 1'b1;
    end
  end

  always @(*) begin
    lineLoader_fire = 1'b0;
    if(io_mem_rsp_valid) begin
      if(when_InstructionCache_l401) begin
        lineLoader_fire = 1'b1;
      end
    end
  end

  always @(*) begin
    io_cpu_prefetch_haltIt = (lineLoader_valid || lineLoader_flushPending);
    if(when_InstructionCache_l338) begin
      io_cpu_prefetch_haltIt = 1'b1;
    end
    if(when_InstructionCache_l342) begin
      io_cpu_prefetch_haltIt = 1'b1;
    end
    if(io_flush) begin
      io_cpu_prefetch_haltIt = 1'b1;
    end
  end

  assign when_InstructionCache_l338 = (! lineLoader_flushCounter[7]);
  assign when_InstructionCache_l342 = (! _zz_when_InstructionCache_l342);
  assign when_InstructionCache_l351 = (lineLoader_flushPending && (! (lineLoader_valid || io_cpu_fetch_isValid)));
  assign io_mem_cmd_fire = (io_mem_cmd_valid && io_mem_cmd_ready);
  assign io_mem_cmd_valid = (lineLoader_valid && (! lineLoader_cmdSent));
  assign io_mem_cmd_payload_address = {lineLoader_address[31 : 5],5'h0};
  assign io_mem_cmd_payload_size = 3'b101;
  assign when_Utils_l515 = (! lineLoader_valid);
  always @(*) begin
    lineLoader_wayToAllocate_willIncrement = 1'b0;
    if(when_Utils_l515) begin
      lineLoader_wayToAllocate_willIncrement = 1'b1;
    end
  end

  assign lineLoader_wayToAllocate_willClear = 1'b0;
  assign lineLoader_wayToAllocate_willOverflowIfInc = 1'b1;
  assign lineLoader_wayToAllocate_willOverflow = (lineLoader_wayToAllocate_willOverflowIfInc && lineLoader_wayToAllocate_willIncrement);
  assign lineLoader_write_tag_0_valid = ((1'b1 && lineLoader_fire) || (! lineLoader_flushCounter[7]));
  assign lineLoader_write_tag_0_payload_address = (lineLoader_flushCounter[7] ? lineLoader_address[11 : 5] : lineLoader_flushCounter[6 : 0]);
  assign lineLoader_write_tag_0_payload_data_valid = lineLoader_flushCounter[7];
  assign lineLoader_write_tag_0_payload_data_error = (lineLoader_hadError || io_mem_rsp_payload_error);
  assign lineLoader_write_tag_0_payload_data_address = lineLoader_address[31 : 12];
  assign lineLoader_write_data_0_valid = (io_mem_rsp_valid && 1'b1);
  assign lineLoader_write_data_0_payload_address = {lineLoader_address[11 : 5],lineLoader_wordIndex};
  assign lineLoader_write_data_0_payload_data = io_mem_rsp_payload_data;
  assign when_InstructionCache_l401 = (lineLoader_wordIndex == 3'b111);
  assign _zz_fetchStage_read_banksValue_0_dataMem = io_cpu_prefetch_pc[11 : 2];
  assign _zz_fetchStage_read_banksValue_0_dataMem_1 = (! io_cpu_fetch_isStuck);
  assign fetchStage_read_banksValue_0_dataMem = _zz_banks_0_port1;
  assign fetchStage_read_banksValue_0_data = fetchStage_read_banksValue_0_dataMem[31 : 0];
  assign _zz_fetchStage_read_waysValues_0_tag_valid = io_cpu_prefetch_pc[11 : 5];
  assign _zz_fetchStage_read_waysValues_0_tag_valid_1 = (! io_cpu_fetch_isStuck);
  assign _zz_fetchStage_read_waysValues_0_tag_valid_2 = _zz_ways_0_tags_port1;
  assign fetchStage_read_waysValues_0_tag_valid = _zz_fetchStage_read_waysValues_0_tag_valid_2[0];
  assign fetchStage_read_waysValues_0_tag_error = _zz_fetchStage_read_waysValues_0_tag_valid_2[1];
  assign fetchStage_read_waysValues_0_tag_address = _zz_fetchStage_read_waysValues_0_tag_valid_2[21 : 2];
  assign fetchStage_hit_hits_0 = (fetchStage_read_waysValues_0_tag_valid && (fetchStage_read_waysValues_0_tag_address == io_cpu_fetch_mmuRsp_physicalAddress[31 : 12]));
  assign fetchStage_hit_valid = (|fetchStage_hit_hits_0);
  assign fetchStage_hit_error = fetchStage_read_waysValues_0_tag_error;
  assign fetchStage_hit_data = fetchStage_read_banksValue_0_data;
  assign fetchStage_hit_word = fetchStage_hit_data;
  assign io_cpu_fetch_data = fetchStage_hit_word;
  assign when_InstructionCache_l435 = (! io_cpu_decode_isStuck);
  assign io_cpu_decode_data = io_cpu_fetch_data_regNextWhen;
  assign io_cpu_fetch_physicalAddress = io_cpu_fetch_mmuRsp_physicalAddress;
  assign when_InstructionCache_l459 = (! io_cpu_decode_isStuck);
  assign when_InstructionCache_l459_1 = (! io_cpu_decode_isStuck);
  assign when_InstructionCache_l459_2 = (! io_cpu_decode_isStuck);
  assign io_cpu_decode_cacheMiss = (! decodeStage_hit_valid);
  assign io_cpu_decode_error = (decodeStage_hit_error || ((! decodeStage_mmuRsp_isPaging) && (decodeStage_mmuRsp_exception || (! decodeStage_mmuRsp_allowExecute))));
  assign io_cpu_decode_mmuRefilling = decodeStage_mmuRsp_refilling;
  assign io_cpu_decode_mmuException = (((! decodeStage_mmuRsp_refilling) && decodeStage_mmuRsp_isPaging) && (decodeStage_mmuRsp_exception || (! decodeStage_mmuRsp_allowExecute)));
  assign io_cpu_decode_physicalAddress = decodeStage_mmuRsp_physicalAddress;
  always @(posedge clk) begin
    if(reset) begin
      lineLoader_valid <= 1'b0;
      lineLoader_hadError <= 1'b0;
      lineLoader_flushPending <= 1'b1;
      lineLoader_cmdSent <= 1'b0;
      lineLoader_wordIndex <= 3'b000;
    end else begin
      if(lineLoader_fire) begin
        lineLoader_valid <= 1'b0;
      end
      if(lineLoader_fire) begin
        lineLoader_hadError <= 1'b0;
      end
      if(io_cpu_fill_valid) begin
        lineLoader_valid <= 1'b1;
      end
      if(io_flush) begin
        lineLoader_flushPending <= 1'b1;
      end
      if(when_InstructionCache_l351) begin
        lineLoader_flushPending <= 1'b0;
      end
      if(io_mem_cmd_fire) begin
        lineLoader_cmdSent <= 1'b1;
      end
      if(lineLoader_fire) begin
        lineLoader_cmdSent <= 1'b0;
      end
      if(io_mem_rsp_valid) begin
        lineLoader_wordIndex <= (lineLoader_wordIndex + 3'b001);
        if(io_mem_rsp_payload_error) begin
          lineLoader_hadError <= 1'b1;
        end
      end
    end
  end

  always @(posedge clk) begin
    if(io_cpu_fill_valid) begin
      lineLoader_address <= io_cpu_fill_payload;
    end
    if(when_InstructionCache_l338) begin
      lineLoader_flushCounter <= (lineLoader_flushCounter + 8'h01);
    end
    _zz_when_InstructionCache_l342 <= lineLoader_flushCounter[7];
    if(when_InstructionCache_l351) begin
      lineLoader_flushCounter <= 8'h0;
    end
    if(when_InstructionCache_l435) begin
      io_cpu_fetch_data_regNextWhen <= io_cpu_fetch_data;
    end
    if(when_InstructionCache_l459) begin
      decodeStage_mmuRsp_physicalAddress <= io_cpu_fetch_mmuRsp_physicalAddress;
      decodeStage_mmuRsp_isIoAccess <= io_cpu_fetch_mmuRsp_isIoAccess;
      decodeStage_mmuRsp_isPaging <= io_cpu_fetch_mmuRsp_isPaging;
      decodeStage_mmuRsp_allowRead <= io_cpu_fetch_mmuRsp_allowRead;
      decodeStage_mmuRsp_allowWrite <= io_cpu_fetch_mmuRsp_allowWrite;
      decodeStage_mmuRsp_allowExecute <= io_cpu_fetch_mmuRsp_allowExecute;
      decodeStage_mmuRsp_exception <= io_cpu_fetch_mmuRsp_exception;
      decodeStage_mmuRsp_refilling <= io_cpu_fetch_mmuRsp_refilling;
      decodeStage_mmuRsp_bypassTranslation <= io_cpu_fetch_mmuRsp_bypassTranslation;
    end
    if(when_InstructionCache_l459_1) begin
      decodeStage_hit_valid <= fetchStage_hit_valid;
    end
    if(when_InstructionCache_l459_2) begin
      decodeStage_hit_error <= fetchStage_hit_error;
    end
  end


endmodule

module PmpSetter (
  input      [31:0]   io_addr,
  output     [24:0]   io_base,
  output     [24:0]   io_mask
);

  wire       [31:0]   _zz_ones;
  wire       [31:0]   ones;

  assign _zz_ones = (io_addr + 32'h00000001);
  assign ones = (io_addr & (~ _zz_ones));
  assign io_base = (io_addr[29 : 5] ^ ones[29 : 5]);
  assign io_mask = (~ {ones[28 : 5],1'b1});

endmodule
